* NGSPICE file created from distance_display.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt distance_display i_clk i_reset i_sensor_echo o_display_anode[0] o_display_anode[1]
+ o_display_anode[2] o_display_anode[3] o_display_cathode[0] o_display_cathode[1]
+ o_display_cathode[2] o_display_cathode[3] o_display_cathode[4] o_display_cathode[5]
+ o_display_cathode[6] o_display_cathode[7] o_io_oeb[0] o_io_oeb[10] o_io_oeb[11]
+ o_io_oeb[12] o_io_oeb[1] o_io_oeb[2] o_io_oeb[3] o_io_oeb[4] o_io_oeb[5] o_io_oeb[6]
+ o_io_oeb[7] o_io_oeb[8] o_io_oeb[9] o_sensor_trigger vccd1 vssd1
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2106_ _2749_/Q _2104_/X _2105_/X vssd1 vssd1 vccd1 vccd1 _2106_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2037_ _2739_/Q vssd1 vssd1 vccd1 vccd1 _2132_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1606_ _1614_/A _1614_/B _1589_/X vssd1 vssd1 vccd1 vccd1 _1606_/X sky130_fd_sc_hd__a21o_1
X_2724_ _2726_/CLK _2724_/D vssd1 vssd1 vccd1 vccd1 _2724_/Q sky130_fd_sc_hd__dfxtp_1
X_2655_ _2809_/Q _2655_/B vssd1 vssd1 vccd1 vccd1 _2655_/X sky130_fd_sc_hd__or2_1
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1468_ _1602_/A vssd1 vssd1 vccd1 vccd1 _1485_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1399_ _1553_/A _1553_/B _1393_/Y vssd1 vssd1 vccd1 vccd1 _1407_/B sky130_fd_sc_hd__a21boi_1
X_1537_ _1684_/A _1523_/Y _1529_/X _1538_/B _1698_/A vssd1 vssd1 vccd1 vccd1 _1537_/X
+ sky130_fd_sc_hd__a311o_1
X_2586_ _2803_/Q _2632_/B _2585_/X _2581_/B vssd1 vssd1 vccd1 vccd1 _2587_/A sky130_fd_sc_hd__a22o_1
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2440_ _2442_/B _2440_/B vssd1 vssd1 vccd1 vccd1 _2441_/A sky130_fd_sc_hd__and2_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2371_ _2699_/Q _2373_/C vssd1 vssd1 vccd1 vccd1 _2699_/D sky130_fd_sc_hd__xor2_1
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2707_ _2807_/CLK _2707_/D vssd1 vssd1 vccd1 vccd1 _2707_/Q sky130_fd_sc_hd__dfxtp_1
X_2638_ _2638_/A vssd1 vssd1 vccd1 vccd1 _2638_/Y sky130_fd_sc_hd__inv_2
X_2569_ _2569_/A _2569_/B vssd1 vssd1 vccd1 vccd1 _2570_/A sky130_fd_sc_hd__and2_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1940_ _2018_/A vssd1 vssd1 vccd1 vccd1 _1940_/Y sky130_fd_sc_hd__inv_2
X_1871_ _1871_/A _1963_/A vssd1 vssd1 vccd1 vccd1 _1871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2423_ _2425_/B _2423_/B vssd1 vssd1 vccd1 vccd1 _2719_/D sky130_fd_sc_hd__nor2_1
X_2285_ _2285_/A vssd1 vssd1 vccd1 vccd1 _2482_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2354_ _2709_/Q _2708_/Q _2711_/Q _2710_/Q vssd1 vssd1 vccd1 vccd1 _2355_/D sky130_fd_sc_hd__or4_1
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2070_ _2146_/A vssd1 vssd1 vccd1 vccd1 _2070_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1923_ _2030_/A _2013_/A vssd1 vssd1 vccd1 vccd1 _1923_/X sky130_fd_sc_hd__or2_1
X_1854_ _1854_/A _1854_/B vssd1 vssd1 vccd1 vccd1 _1854_/Y sky130_fd_sc_hd__nor2_1
X_1785_ _1779_/Y _1812_/S _1784_/X vssd1 vssd1 vccd1 vccd1 _1807_/B sky130_fd_sc_hd__o21ai_2
X_2406_ _2712_/Q _2407_/C vssd1 vssd1 vccd1 vccd1 _2712_/D sky130_fd_sc_hd__xor2_1
X_2337_ _2688_/Q _2342_/C vssd1 vssd1 vccd1 vccd1 _2339_/A sky130_fd_sc_hd__or2_1
X_2268_ _2674_/Q _2673_/Q vssd1 vssd1 vccd1 vccd1 _2270_/C sky130_fd_sc_hd__nand2_1
X_2199_ _2657_/Q _2658_/Q vssd1 vssd1 vccd1 vccd1 _2199_/Y sky130_fd_sc_hd__nor2_4
XFILLER_40_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1570_ _1570_/A _1570_/B vssd1 vssd1 vccd1 vccd1 _1573_/A sky130_fd_sc_hd__nor2_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _2146_/A vssd1 vssd1 vccd1 vccd1 _2122_/X sky130_fd_sc_hd__clkbuf_2
X_2053_ _2053_/A _2154_/A vssd1 vssd1 vccd1 vccd1 _2149_/B sky130_fd_sc_hd__and2_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1768_ _1791_/B _1766_/X _1767_/X vssd1 vssd1 vccd1 vccd1 _1768_/Y sky130_fd_sc_hd__a21oi_1
X_1906_ _1890_/A _1889_/X _1905_/Y _1985_/A vssd1 vssd1 vccd1 vccd1 _1906_/X sky130_fd_sc_hd__o211a_1
X_1837_ _2053_/A _1837_/B vssd1 vssd1 vccd1 vccd1 _1857_/A sky130_fd_sc_hd__xnor2_2
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1699_ _1699_/A _1699_/B vssd1 vssd1 vccd1 vccd1 _1721_/S sky130_fd_sc_hd__xnor2_2
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput7 _2223_/X vssd1 vssd1 vccd1 vccd1 o_display_cathode[1] sky130_fd_sc_hd__buf_2
XFILLER_56_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1622_ _1624_/B _1624_/C _1899_/B vssd1 vssd1 vccd1 vccd1 _1641_/A sky130_fd_sc_hd__a21oi_2
X_2671_ _2727_/CLK _2671_/D vssd1 vssd1 vccd1 vccd1 _2671_/Q sky130_fd_sc_hd__dfxtp_1
X_2740_ _2759_/CLK _2740_/D _2459_/Y vssd1 vssd1 vccd1 vccd1 _2740_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1484_ _1485_/B _1602_/B _1485_/A vssd1 vssd1 vccd1 vccd1 _1489_/A sky130_fd_sc_hd__a21o_1
X_1553_ _1553_/A _1553_/B vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__nand2_2
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2105_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2105_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2036_ _2036_/A vssd1 vssd1 vccd1 vccd1 _2761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2723_ _2726_/CLK _2723_/D vssd1 vssd1 vccd1 vccd1 _2723_/Q sky130_fd_sc_hd__dfxtp_1
X_1605_ _1899_/A _1599_/X _1612_/B vssd1 vssd1 vccd1 vccd1 _1608_/A sky130_fd_sc_hd__o21ai_1
X_1536_ _2741_/Q _1536_/B vssd1 vssd1 vccd1 vccd1 _1698_/A sky130_fd_sc_hd__xnor2_1
X_2585_ _2799_/Q _2807_/Q _2787_/Q vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__mux2_1
X_2654_ _2808_/Q _2249_/A _2653_/X _2244_/A vssd1 vssd1 vccd1 vccd1 _2654_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1467_ _1590_/A _1467_/B vssd1 vssd1 vccd1 vccd1 _1602_/A sky130_fd_sc_hd__or2_1
X_1398_ _1391_/Y _1396_/Y _1553_/A vssd1 vssd1 vccd1 vccd1 _1412_/A sky130_fd_sc_hd__o21a_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2019_ _2765_/Q _2018_/Y _2032_/S vssd1 vssd1 vccd1 vccd1 _2020_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2370_ _2370_/A _2373_/C vssd1 vssd1 vccd1 vccd1 _2698_/D sky130_fd_sc_hd__nor2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2706_ _2757_/CLK _2706_/D vssd1 vssd1 vccd1 vccd1 _2706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1519_ _1519_/A _1524_/A vssd1 vssd1 vccd1 vccd1 _1520_/S sky130_fd_sc_hd__xnor2_1
X_2499_ _2774_/Q _2779_/Q _2778_/Q vssd1 vssd1 vccd1 vccd1 _2502_/B sky130_fd_sc_hd__and3_1
X_2637_ _2804_/Q _2617_/X _2635_/X _2636_/X vssd1 vssd1 vccd1 vccd1 _2804_/D sky130_fd_sc_hd__o211a_1
X_2568_ _2796_/Q _2567_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2569_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1870_ _1870_/A _1870_/B vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2422_ _2718_/Q _2421_/C _2719_/Q vssd1 vssd1 vccd1 vccd1 _2423_/B sky130_fd_sc_hd__a21oi_1
X_2353_ _2705_/Q _2704_/Q _2707_/Q _2706_/Q vssd1 vssd1 vccd1 vccd1 _2355_/C sky130_fd_sc_hd__or4_1
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2284_ _2666_/Q _2667_/Q _2284_/C vssd1 vssd1 vccd1 vccd1 _2288_/B sky130_fd_sc_hd__and3_1
XFILLER_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1999_ _1940_/Y _2022_/A _2026_/A _2025_/B _2025_/A vssd1 vssd1 vccd1 vccd1 _2013_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1922_ _1935_/C vssd1 vssd1 vccd1 vccd1 _2013_/A sky130_fd_sc_hd__clkbuf_2
X_1853_ _1862_/A _1853_/B vssd1 vssd1 vccd1 vccd1 _1856_/A sky130_fd_sc_hd__nor2_1
X_1784_ _1754_/X _1755_/Y _1783_/Y vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__a21o_1
X_2336_ _2336_/A _2342_/C vssd1 vssd1 vccd1 vccd1 _2687_/D sky130_fd_sc_hd__nor2_1
X_2405_ _2407_/C _2405_/B vssd1 vssd1 vccd1 vccd1 _2711_/D sky130_fd_sc_hd__nor2_1
X_2267_ _2680_/Q _2679_/Q _2682_/Q _2681_/Q vssd1 vssd1 vccd1 vccd1 _2271_/C sky130_fd_sc_hd__or4_1
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2198_ _2198_/A vssd1 vssd1 vccd1 vccd1 _2775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2121_ _2121_/A _2121_/B vssd1 vssd1 vccd1 vccd1 _2121_/X sky130_fd_sc_hd__or2_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2052_ _2052_/A _2052_/B _2159_/A vssd1 vssd1 vccd1 vccd1 _2154_/A sky130_fd_sc_hd__and3_1
X_1905_ _1948_/A _1963_/A _1976_/A _1905_/D vssd1 vssd1 vccd1 vccd1 _1905_/Y sky130_fd_sc_hd__nor4_1
X_1698_ _1698_/A _1902_/B vssd1 vssd1 vccd1 vccd1 _1699_/B sky130_fd_sc_hd__or2b_1
X_1767_ _1767_/A _1767_/B _1767_/C _1792_/A vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__and4_1
X_1836_ _1887_/A _2052_/A _1834_/B vssd1 vssd1 vccd1 vccd1 _1837_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2319_ _2319_/A _2321_/B vssd1 vssd1 vccd1 vccd1 _2680_/D sky130_fd_sc_hd__nor2_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2820__23 vssd1 vssd1 vccd1 vccd1 _2820__23/HI o_io_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput8 _2226_/X vssd1 vssd1 vccd1 vccd1 o_display_cathode[2] sky130_fd_sc_hd__buf_2
Xoutput10 _2231_/Y vssd1 vssd1 vccd1 vccd1 o_display_cathode[4] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_i_clk clkbuf_3_7_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _2673_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1621_ _1589_/X _1594_/X _1618_/X _1620_/Y vssd1 vssd1 vccd1 vccd1 _1624_/C sky130_fd_sc_hd__a2bb2o_2
X_1552_ _1552_/A vssd1 vssd1 vccd1 vccd1 _1561_/A sky130_fd_sc_hd__inv_2
X_2670_ _2727_/CLK _2670_/D vssd1 vssd1 vccd1 vccd1 _2670_/Q sky130_fd_sc_hd__dfxtp_1
X_1483_ _1483_/A _1483_/B _1546_/B vssd1 vssd1 vccd1 vccd1 _1496_/B sky130_fd_sc_hd__and3_1
X_2104_ _2104_/A _2110_/A vssd1 vssd1 vccd1 vccd1 _2104_/X sky130_fd_sc_hd__and2_1
XFILLER_39_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2035_ _2761_/Q _2034_/Y _2695_/Q vssd1 vssd1 vccd1 vccd1 _2036_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2799_ _2806_/CLK _2799_/D vssd1 vssd1 vccd1 vccd1 _2799_/Q sky130_fd_sc_hd__dfxtp_1
X_1819_ _1818_/X _1817_/Y _1819_/S vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2722_ _2726_/CLK _2722_/D vssd1 vssd1 vccd1 vccd1 _2722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1604_ _1612_/A _1604_/B vssd1 vssd1 vccd1 vccd1 _1604_/Y sky130_fd_sc_hd__xnor2_1
X_1535_ _1749_/A _2056_/A _1695_/B vssd1 vssd1 vccd1 vccd1 _1536_/B sky130_fd_sc_hd__a21oi_1
X_2653_ _2525_/A _2183_/A _2638_/Y _2183_/Y _2809_/Q vssd1 vssd1 vccd1 vccd1 _2653_/X
+ sky130_fd_sc_hd__a32o_1
X_2584_ _2800_/Q _2580_/Y _2583_/X vssd1 vssd1 vccd1 vccd1 _2610_/A sky130_fd_sc_hd__a21oi_1
X_1466_ _1462_/Y _1590_/B _1458_/X _1457_/Y vssd1 vssd1 vccd1 vccd1 _1467_/B sky130_fd_sc_hd__a211oi_1
X_1397_ _1403_/A _1393_/Y _1391_/A _1391_/B vssd1 vssd1 vccd1 vccd1 _1553_/A sky130_fd_sc_hd__a22o_1
X_2018_ _2018_/A _2018_/B vssd1 vssd1 vccd1 vccd1 _2018_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_12_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2705_ _2807_/CLK _2705_/D vssd1 vssd1 vccd1 vccd1 _2705_/Q sky130_fd_sc_hd__dfxtp_1
X_2636_ _2636_/A vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__clkbuf_2
X_1449_ _1571_/A _1571_/B _1447_/A _1444_/A vssd1 vssd1 vccd1 vccd1 _1449_/X sky130_fd_sc_hd__o2bb2a_1
X_1518_ _1518_/A _1518_/B vssd1 vssd1 vccd1 vccd1 _1518_/Y sky130_fd_sc_hd__nand2_1
X_2498_ _2778_/Q _2186_/X _2497_/Y vssd1 vssd1 vccd1 vccd1 _2778_/D sky130_fd_sc_hd__o21a_1
X_2567_ _2768_/Q _2795_/Q _2598_/A vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2283_ _2283_/A _2283_/B vssd1 vssd1 vccd1 vccd1 _2666_/D sky130_fd_sc_hd__nor2_1
X_2421_ _2719_/Q _2718_/Q _2421_/C vssd1 vssd1 vccd1 vccd1 _2425_/B sky130_fd_sc_hd__and3_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2352_ _2697_/Q _2696_/D _2699_/Q _2698_/Q vssd1 vssd1 vccd1 vccd1 _2355_/B sky130_fd_sc_hd__or4_1
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2619_ _2801_/Q _2576_/X _2577_/X _2598_/X _2800_/Q vssd1 vssd1 vccd1 vccd1 _2623_/B
+ sky130_fd_sc_hd__a32o_1
X_1998_ _1909_/X _1923_/X _1996_/Y _1997_/Y vssd1 vssd1 vccd1 vccd1 _1998_/X sky130_fd_sc_hd__a31o_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1921_ _1936_/A _1924_/A _1930_/A _1930_/B _1920_/Y vssd1 vssd1 vccd1 vccd1 _1935_/C
+ sky130_fd_sc_hd__o41a_1
X_1852_ _1852_/A _1852_/B vssd1 vssd1 vccd1 vccd1 _1853_/B sky130_fd_sc_hd__xnor2_1
X_1783_ _1758_/X _1754_/X _1755_/Y vssd1 vssd1 vccd1 vccd1 _1783_/Y sky130_fd_sc_hd__a21oi_1
X_2335_ _2687_/Q _2335_/B vssd1 vssd1 vccd1 vccd1 _2342_/C sky130_fd_sc_hd__and2_1
X_2266_ _2684_/Q _2683_/Q _2686_/Q _2685_/Q vssd1 vssd1 vccd1 vccd1 _2271_/B sky130_fd_sc_hd__or4_1
X_2404_ _2711_/Q _2404_/B vssd1 vssd1 vccd1 vccd1 _2405_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2197_ _2546_/A _2197_/B vssd1 vssd1 vccd1 vccd1 _2198_/A sky130_fd_sc_hd__and2_1
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_11_0_i_clk clkbuf_3_5_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _2727_/CLK sky130_fd_sc_hd__clkbuf_2
X_2120_ _2121_/A _2121_/B vssd1 vssd1 vccd1 vccd1 _2120_/Y sky130_fd_sc_hd__nand2_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ _2731_/Q _2730_/Q _2165_/A vssd1 vssd1 vccd1 vccd1 _2159_/A sky130_fd_sc_hd__and3_1
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1904_ _1904_/A _1917_/A _1928_/A _1904_/D vssd1 vssd1 vccd1 vccd1 _1905_/D sky130_fd_sc_hd__or4_1
X_1835_ _2734_/Q vssd1 vssd1 vccd1 vccd1 _2053_/A sky130_fd_sc_hd__clkbuf_2
X_1697_ _1684_/A _1523_/Y _1529_/X _1538_/B vssd1 vssd1 vccd1 vccd1 _1699_/A sky130_fd_sc_hd__a31o_1
X_1766_ _1766_/A _1766_/B vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__or2_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2318_ _2680_/Q _2679_/Q _2318_/C vssd1 vssd1 vccd1 vccd1 _2321_/B sky130_fd_sc_hd__and3_1
X_2249_ _2249_/A _2636_/A vssd1 vssd1 vccd1 vccd1 _2250_/A sky130_fd_sc_hd__and2_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput11 _2232_/X vssd1 vssd1 vccd1 vccd1 o_display_cathode[5] sky130_fd_sc_hd__buf_2
Xoutput9 _2229_/X vssd1 vssd1 vccd1 vccd1 o_display_cathode[3] sky130_fd_sc_hd__buf_2
XFILLER_0_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1620_ _1620_/A _1620_/B vssd1 vssd1 vccd1 vccd1 _1620_/Y sky130_fd_sc_hd__xnor2_1
X_1551_ _1551_/A _1551_/B vssd1 vssd1 vccd1 vccd1 _1552_/A sky130_fd_sc_hd__nand2_1
X_1482_ _1485_/C _1480_/X _1602_/B vssd1 vssd1 vccd1 vccd1 _1546_/B sky130_fd_sc_hd__a21bo_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2103_ _2088_/X _2101_/Y _2102_/X _2099_/X _2102_/A vssd1 vssd1 vccd1 vccd1 _2750_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2034_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2034_/Y sky130_fd_sc_hd__inv_2
X_2798_ _2807_/CLK _2798_/D vssd1 vssd1 vccd1 vccd1 _2798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1818_ _1817_/Y _1818_/B vssd1 vssd1 vccd1 vccd1 _1818_/X sky130_fd_sc_hd__and2b_1
X_1749_ _1749_/A vssd1 vssd1 vccd1 vccd1 _1823_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2721_ _2806_/CLK _2721_/D vssd1 vssd1 vccd1 vccd1 _2721_/Q sky130_fd_sc_hd__dfxtp_1
X_2652_ _2808_/Q _2655_/B _2651_/X _2636_/X vssd1 vssd1 vccd1 vccd1 _2808_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1603_ _1899_/B vssd1 vssd1 vccd1 vccd1 _1603_/Y sky130_fd_sc_hd__inv_2
X_1465_ _1470_/C vssd1 vssd1 vccd1 vccd1 _1590_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1534_ _1805_/B _1511_/D _1749_/A vssd1 vssd1 vccd1 vccd1 _1695_/B sky130_fd_sc_hd__o21a_1
X_2583_ _2808_/Q _2195_/X _2629_/S _2804_/Q vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__a22o_1
X_1396_ _1403_/A _1393_/Y _1553_/B vssd1 vssd1 vccd1 vccd1 _1396_/Y sky130_fd_sc_hd__a21oi_1
X_2017_ _2022_/A _2026_/A _2025_/B _2025_/A vssd1 vssd1 vccd1 vccd1 _2018_/B sky130_fd_sc_hd__o31a_1
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2704_ _2807_/CLK _2704_/D vssd1 vssd1 vccd1 vccd1 _2704_/Q sky130_fd_sc_hd__dfxtp_1
X_2635_ _2803_/Q _2248_/A _2634_/X _2244_/A _2625_/X vssd1 vssd1 vccd1 vccd1 _2635_/X
+ sky130_fd_sc_hd__a221o_1
X_1448_ _1448_/A _1448_/B vssd1 vssd1 vccd1 vccd1 _1448_/X sky130_fd_sc_hd__and2_1
X_1517_ _1499_/Y _1516_/X _1545_/A vssd1 vssd1 vccd1 vccd1 _1518_/B sky130_fd_sc_hd__a21boi_1
X_2497_ _2503_/A _2497_/B vssd1 vssd1 vccd1 vccd1 _2497_/Y sky130_fd_sc_hd__nor2_1
X_2566_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2795_/D sky130_fd_sc_hd__clkbuf_1
X_1379_ _2754_/Q vssd1 vssd1 vccd1 vccd1 _2064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2420_ _2718_/Q _2421_/C vssd1 vssd1 vccd1 vccd1 _2718_/D sky130_fd_sc_hd__xor2_1
X_2282_ _2666_/Q _2284_/C vssd1 vssd1 vccd1 vccd1 _2283_/B sky130_fd_sc_hd__nor2_1
X_2351_ _2696_/Q vssd1 vssd1 vccd1 vccd1 _2696_/D sky130_fd_sc_hd__inv_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1997_ _2001_/A vssd1 vssd1 vccd1 vccd1 _1997_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2618_ _2618_/A vssd1 vssd1 vccd1 vccd1 _2625_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2549_ _2764_/Q _2791_/Q _2553_/S vssd1 vssd1 vccd1 vccd1 _2549_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1920_ _1920_/A _1920_/B vssd1 vssd1 vccd1 vccd1 _1920_/Y sky130_fd_sc_hd__xnor2_1
X_1851_ _1851_/A _1928_/A vssd1 vssd1 vccd1 vccd1 _1852_/B sky130_fd_sc_hd__nand2_1
X_2403_ _2711_/Q _2404_/B vssd1 vssd1 vccd1 vccd1 _2407_/C sky130_fd_sc_hd__and2_1
X_1782_ _1758_/X _1780_/Y _1776_/A _1781_/Y vssd1 vssd1 vccd1 vccd1 _1812_/S sky130_fd_sc_hd__a31oi_2
X_2265_ _2688_/Q _2687_/Q _2690_/Q _2689_/Q vssd1 vssd1 vccd1 vccd1 _2271_/A sky130_fd_sc_hd__or4_1
X_2334_ _2687_/Q _2335_/B vssd1 vssd1 vccd1 vccd1 _2336_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2196_ _2771_/Q _2772_/Q _2195_/X _2773_/Q vssd1 vssd1 vccd1 vccd1 _2197_/B sky130_fd_sc_hd__a22o_1
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ _2735_/Q vssd1 vssd1 vccd1 vccd1 _2149_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1765_ _1764_/B _1764_/C _1767_/A vssd1 vssd1 vccd1 vccd1 _1766_/B sky130_fd_sc_hd__a21oi_1
X_1834_ _2052_/A _1834_/B vssd1 vssd1 vccd1 vccd1 _1870_/B sky130_fd_sc_hd__xnor2_2
X_1903_ _1903_/A _1903_/B _1903_/C vssd1 vssd1 vccd1 vccd1 _1904_/D sky130_fd_sc_hd__or3_1
X_1696_ _1696_/A _1722_/A vssd1 vssd1 vccd1 vccd1 _1720_/A sky130_fd_sc_hd__or2b_1
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2317_ _2679_/Q _2318_/C _2680_/Q vssd1 vssd1 vccd1 vccd1 _2319_/A sky130_fd_sc_hd__a21oi_1
X_2248_ _2248_/A vssd1 vssd1 vccd1 vccd1 _2249_/A sky130_fd_sc_hd__clkbuf_2
X_2179_ _2788_/Q vssd1 vssd1 vccd1 vccd1 _2632_/A sky130_fd_sc_hd__inv_2
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput12 _2233_/Y vssd1 vssd1 vccd1 vccd1 o_display_cathode[6] sky130_fd_sc_hd__buf_2
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2811__14 vssd1 vssd1 vccd1 vccd1 _2811__14/HI o_io_oeb[0] sky130_fd_sc_hd__conb_1
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1550_ _1563_/A vssd1 vssd1 vccd1 vccd1 _1578_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1481_ _1352_/A _1471_/A _1471_/B _1477_/A _1477_/B vssd1 vssd1 vccd1 vccd1 _1602_/B
+ sky130_fd_sc_hd__a311o_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2102_ _2102_/A _2102_/B vssd1 vssd1 vccd1 vccd1 _2102_/X sky130_fd_sc_hd__or2_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_i_clk clkbuf_4_9_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2807_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1748_ _2738_/Q vssd1 vssd1 vccd1 vccd1 _2055_/A sky130_fd_sc_hd__clkbuf_2
X_2797_ _2802_/CLK _2797_/D vssd1 vssd1 vccd1 vccd1 _2797_/Q sky130_fd_sc_hd__dfxtp_1
X_1817_ _1910_/A _1817_/B _1920_/A vssd1 vssd1 vccd1 vccd1 _1817_/Y sky130_fd_sc_hd__nand3_1
X_1679_ _1901_/B _1679_/B vssd1 vssd1 vccd1 vccd1 _1680_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1602_ _1602_/A _1602_/B vssd1 vssd1 vccd1 vccd1 _1899_/B sky130_fd_sc_hd__nand2_2
X_2720_ _2806_/CLK _2720_/D vssd1 vssd1 vccd1 vccd1 _2720_/Q sky130_fd_sc_hd__dfxtp_1
X_2651_ _2807_/Q _2248_/A _2650_/X _2242_/A _2625_/A vssd1 vssd1 vccd1 vccd1 _2651_/X
+ sky130_fd_sc_hd__a221o_1
X_2582_ _2590_/A _2582_/B vssd1 vssd1 vccd1 vccd1 _2629_/S sky130_fd_sc_hd__nor2_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1464_ _1445_/X _1447_/X _1463_/Y vssd1 vssd1 vccd1 vccd1 _1470_/C sky130_fd_sc_hd__a21oi_1
X_1395_ _1394_/Y _1394_/B _1395_/S vssd1 vssd1 vccd1 vccd1 _1553_/B sky130_fd_sc_hd__mux2_1
X_1533_ _2740_/Q vssd1 vssd1 vccd1 vccd1 _2056_/A sky130_fd_sc_hd__clkbuf_2
X_2016_ _2016_/A vssd1 vssd1 vccd1 vccd1 _2766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1516_ _1504_/A _1519_/A _1545_/B vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__a21o_1
X_2703_ _2807_/CLK _2703_/D vssd1 vssd1 vccd1 vccd1 _2703_/Q sky130_fd_sc_hd__dfxtp_1
X_2565_ _2569_/A _2565_/B vssd1 vssd1 vccd1 vccd1 _2566_/A sky130_fd_sc_hd__and2_1
X_2634_ _2804_/Q _2632_/Y _2633_/Y _2521_/X vssd1 vssd1 vccd1 vccd1 _2634_/X sky130_fd_sc_hd__a22o_1
X_1447_ _1447_/A _1456_/A vssd1 vssd1 vccd1 vccd1 _1447_/X sky130_fd_sc_hd__xor2_1
X_1378_ _1378_/A _1549_/A _1549_/B vssd1 vssd1 vccd1 vccd1 _1383_/C sky130_fd_sc_hd__and3_1
XFILLER_4_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2496_ _2774_/Q _2778_/Q vssd1 vssd1 vccd1 vccd1 _2497_/B sky130_fd_sc_hd__and2_1
Xclkbuf_3_6_0_i_clk clkbuf_3_7_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_i_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2281_ _2666_/Q _2284_/C vssd1 vssd1 vccd1 vccd1 _2283_/A sky130_fd_sc_hd__and2_1
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2350_ _2703_/Q _2702_/Q _2701_/Q _2700_/Q vssd1 vssd1 vccd1 vccd1 _2355_/A sky130_fd_sc_hd__or4bb_1
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1996_ _1940_/Y _2022_/A _2026_/A _2025_/B _2025_/A vssd1 vssd1 vccd1 vccd1 _1996_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2617_ _2655_/B vssd1 vssd1 vccd1 vccd1 _2617_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2548_ _2571_/A vssd1 vssd1 vccd1 vccd1 _2569_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2479_ _2481_/A vssd1 vssd1 vccd1 vccd1 _2479_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1850_ _1850_/A vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__clkbuf_2
X_1781_ _1776_/A _1903_/B _1780_/Y vssd1 vssd1 vccd1 vccd1 _1781_/Y sky130_fd_sc_hd__a21oi_1
X_2333_ _2333_/A _2335_/B vssd1 vssd1 vccd1 vccd1 _2686_/D sky130_fd_sc_hd__nor2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2402_ _2404_/B _2402_/B vssd1 vssd1 vccd1 vccd1 _2710_/D sky130_fd_sc_hd__nor2_1
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2817__20 vssd1 vssd1 vccd1 vccd1 _2817__20/HI o_io_oeb[6] sky130_fd_sc_hd__conb_1
X_2264_ _2676_/Q _2675_/Q _2678_/Q _2677_/Q vssd1 vssd1 vccd1 vccd1 _2272_/C sky130_fd_sc_hd__or4_1
X_2195_ _2632_/A _2581_/A _2581_/B vssd1 vssd1 vccd1 vccd1 _2195_/X sky130_fd_sc_hd__and3_1
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1979_ _1978_/A _1978_/C _1978_/B vssd1 vssd1 vccd1 vccd1 _1979_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_i_clk clkbuf_2_3_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1902_ _1902_/A _1902_/B _1731_/A _1901_/X vssd1 vssd1 vccd1 vccd1 _1903_/C sky130_fd_sc_hd__or4bb_1
X_1764_ _1767_/A _1764_/B _1764_/C vssd1 vssd1 vccd1 vccd1 _1766_/A sky130_fd_sc_hd__and3_1
X_1833_ _2733_/Q vssd1 vssd1 vccd1 vccd1 _2052_/A sky130_fd_sc_hd__clkbuf_2
X_2316_ _2679_/Q _2318_/C vssd1 vssd1 vccd1 vccd1 _2679_/D sky130_fd_sc_hd__xor2_1
X_1695_ _2056_/A _1695_/B vssd1 vssd1 vccd1 vccd1 _1722_/A sky130_fd_sc_hd__xnor2_2
Xclkbuf_4_5_0_i_clk clkbuf_4_5_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2769_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2247_ _2553_/S vssd1 vssd1 vccd1 vccd1 _2248_/A sky130_fd_sc_hd__clkbuf_2
X_2178_ _2581_/B vssd1 vssd1 vccd1 vccd1 _2183_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput13 _2770_/Q vssd1 vssd1 vccd1 vccd1 o_sensor_trigger sky130_fd_sc_hd__buf_2
XFILLER_0_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1480_ _1352_/A _1471_/X _1485_/B vssd1 vssd1 vccd1 vccd1 _1480_/X sky130_fd_sc_hd__a21o_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2101_ _2102_/A _2102_/B vssd1 vssd1 vccd1 vccd1 _2101_/Y sky130_fd_sc_hd__nand2_1
X_2032_ _2762_/Q _2031_/Y _2032_/S vssd1 vssd1 vccd1 vccd1 _2033_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1678_ _1685_/A _1902_/A vssd1 vssd1 vccd1 vccd1 _1688_/A sky130_fd_sc_hd__or2_1
X_1747_ _1744_/A _1758_/A _1746_/Y vssd1 vssd1 vccd1 vccd1 _1755_/B sky130_fd_sc_hd__a21oi_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1816_ _1917_/A _1918_/A vssd1 vssd1 vccd1 vccd1 _1912_/A sky130_fd_sc_hd__or2_2
X_2796_ _2805_/CLK _2796_/D vssd1 vssd1 vccd1 vccd1 _2796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_i_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1601_ _1899_/A _1604_/B vssd1 vssd1 vccd1 vccd1 _1626_/B sky130_fd_sc_hd__xnor2_2
X_1532_ _1684_/A _1684_/B _1523_/Y vssd1 vssd1 vccd1 vccd1 _1538_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_0_0_i_clk clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
X_2581_ _2581_/A _2581_/B vssd1 vssd1 vccd1 vccd1 _2582_/B sky130_fd_sc_hd__or2_1
X_2650_ _2525_/A _2183_/A _2633_/Y _2183_/Y _2808_/Q vssd1 vssd1 vccd1 vccd1 _2650_/X
+ sky130_fd_sc_hd__a32o_1
X_1463_ _1450_/X _1445_/X _1447_/X vssd1 vssd1 vccd1 vccd1 _1463_/Y sky130_fd_sc_hd__a21oi_1
X_1394_ _1394_/A _1394_/B vssd1 vssd1 vccd1 vccd1 _1394_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2015_ _2766_/Q _2013_/Y _2032_/S vssd1 vssd1 vccd1 vccd1 _2016_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2779_ _2783_/CLK _2779_/D vssd1 vssd1 vccd1 vccd1 _2779_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_2_0_i_clk clkbuf_3_3_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2702_ _2807_/CLK _2702_/D vssd1 vssd1 vccd1 vccd1 _2702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1515_ _1524_/A _1524_/B _1530_/A vssd1 vssd1 vccd1 vccd1 _1518_/A sky130_fd_sc_hd__or3_1
X_2633_ _2633_/A vssd1 vssd1 vccd1 vccd1 _2633_/Y sky130_fd_sc_hd__inv_2
X_2495_ _2511_/A vssd1 vssd1 vccd1 vccd1 _2495_/Y sky130_fd_sc_hd__inv_2
X_2564_ _2795_/Q _2563_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2565_/B sky130_fd_sc_hd__mux2_1
X_1446_ _1446_/A _1446_/B vssd1 vssd1 vccd1 vccd1 _1447_/A sky130_fd_sc_hd__or2_1
X_1377_ _1549_/A _1549_/B _1378_/A vssd1 vssd1 vccd1 vccd1 _1383_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2280_ _2280_/A vssd1 vssd1 vccd1 vccd1 _2665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2616_ _2616_/A vssd1 vssd1 vccd1 vccd1 _2800_/D sky130_fd_sc_hd__clkbuf_1
X_1995_ _1995_/A vssd1 vssd1 vccd1 vccd1 _2025_/A sky130_fd_sc_hd__clkinv_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1429_ _1435_/A _1557_/C _1440_/A vssd1 vssd1 vccd1 vccd1 _1446_/A sky130_fd_sc_hd__a21oi_1
X_2478_ _2481_/A vssd1 vssd1 vccd1 vccd1 _2478_/Y sky130_fd_sc_hd__inv_2
X_2547_ _2547_/A vssd1 vssd1 vccd1 vccd1 _2791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1780_ _1744_/A _1746_/Y _1728_/X _1755_/B vssd1 vssd1 vccd1 vccd1 _1780_/Y sky130_fd_sc_hd__a31oi_2
X_2332_ _2686_/Q _2685_/Q _2332_/C vssd1 vssd1 vccd1 vccd1 _2335_/B sky130_fd_sc_hd__and3_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2401_ _2709_/Q _2400_/C _2710_/Q vssd1 vssd1 vccd1 vccd1 _2402_/B sky130_fd_sc_hd__a21oi_1
X_2263_ _2670_/Q _2669_/Q _2672_/Q _2671_/Q vssd1 vssd1 vccd1 vccd1 _2272_/B sky130_fd_sc_hd__or4_1
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2194_ _2571_/A vssd1 vssd1 vccd1 vccd1 _2546_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_i_clk clkbuf_4_1_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2793_/CLK sky130_fd_sc_hd__clkbuf_2
X_1978_ _1978_/A _1978_/B _1978_/C vssd1 vssd1 vccd1 vccd1 _1978_/Y sky130_fd_sc_hd__nand3_1
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1901_ _1901_/A _1901_/B _1901_/C vssd1 vssd1 vccd1 vccd1 _1901_/X sky130_fd_sc_hd__and3_1
X_1832_ _1834_/B _1829_/Y _2041_/A _1831_/Y vssd1 vssd1 vccd1 vccd1 _1877_/A sky130_fd_sc_hd__o2bb2a_1
X_1694_ _1698_/A _1902_/B vssd1 vssd1 vccd1 vccd1 _1696_/A sky130_fd_sc_hd__xor2_1
X_1763_ _1767_/B _1767_/C _1792_/A _1763_/D vssd1 vssd1 vccd1 vccd1 _1791_/B sky130_fd_sc_hd__nand4_1
X_2315_ _2315_/A _2318_/C vssd1 vssd1 vccd1 vccd1 _2678_/D sky130_fd_sc_hd__nor2_1
X_2246_ _2775_/Q vssd1 vssd1 vccd1 vccd1 _2553_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2177_ _2786_/Q vssd1 vssd1 vccd1 vccd1 _2581_/B sky130_fd_sc_hd__inv_2
XFILLER_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2100_ _2088_/X _2097_/Y _2098_/X _2099_/X _2751_/Q vssd1 vssd1 vccd1 vccd1 _2751_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2031_ _2031_/A _2031_/B vssd1 vssd1 vccd1 vccd1 _2031_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1815_ _1904_/A _2006_/A vssd1 vssd1 vccd1 vccd1 _1918_/A sky130_fd_sc_hd__xnor2_1
X_2795_ _2805_/CLK _2795_/D vssd1 vssd1 vccd1 vccd1 _2795_/Q sky130_fd_sc_hd__dfxtp_1
X_1677_ _1677_/A _1684_/B vssd1 vssd1 vccd1 vccd1 _1902_/A sky130_fd_sc_hd__nand2_1
X_1746_ _1756_/B vssd1 vssd1 vccd1 vccd1 _1746_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2229_ _2229_/A vssd1 vssd1 vccd1 vccd1 _2229_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1600_ _1589_/X _1594_/X _1599_/X vssd1 vssd1 vccd1 vccd1 _1604_/B sky130_fd_sc_hd__o21a_1
X_1462_ _1462_/A _1470_/A vssd1 vssd1 vccd1 vccd1 _1462_/Y sky130_fd_sc_hd__nand2_1
X_1531_ _1539_/A _1539_/B _1529_/A _1529_/B vssd1 vssd1 vccd1 vccd1 _1684_/B sky130_fd_sc_hd__a211o_1
X_2580_ _2590_/A _2581_/A _2786_/Q vssd1 vssd1 vccd1 vccd1 _2580_/Y sky130_fd_sc_hd__nor3_1
X_1393_ _2064_/A _1393_/B vssd1 vssd1 vccd1 vccd1 _1393_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2014_ _2695_/Q vssd1 vssd1 vccd1 vccd1 _2032_/S sky130_fd_sc_hd__clkbuf_2
X_2778_ _2783_/CLK _2778_/D vssd1 vssd1 vccd1 vccd1 _2778_/Q sky130_fd_sc_hd__dfxtp_1
X_1729_ _1756_/A _1756_/B _1728_/X vssd1 vssd1 vccd1 vccd1 _1758_/A sky130_fd_sc_hd__a21o_1
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2701_ _2806_/CLK _2701_/D vssd1 vssd1 vccd1 vccd1 _2701_/Q sky130_fd_sc_hd__dfxtp_1
X_2632_ _2632_/A _2632_/B vssd1 vssd1 vccd1 vccd1 _2632_/Y sky130_fd_sc_hd__nand2_1
X_1445_ _1474_/A _1456_/A _1456_/B vssd1 vssd1 vccd1 vccd1 _1445_/X sky130_fd_sc_hd__or3_1
X_1514_ _2058_/A _1514_/B vssd1 vssd1 vccd1 vccd1 _1530_/A sky130_fd_sc_hd__xnor2_2
X_2563_ _2767_/Q _2794_/Q _2598_/A vssd1 vssd1 vccd1 vccd1 _2563_/X sky130_fd_sc_hd__mux2_1
X_2494_ _2494_/A vssd1 vssd1 vccd1 vccd1 _2494_/Y sky130_fd_sc_hd__inv_2
X_1376_ _2756_/Q _1376_/B vssd1 vssd1 vccd1 vccd1 _1378_/A sky130_fd_sc_hd__xor2_1
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ _2031_/A _2029_/A _2029_/B vssd1 vssd1 vccd1 vccd1 _2025_/B sky130_fd_sc_hd__or3_2
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2615_ _2645_/A _2615_/B vssd1 vssd1 vccd1 vccd1 _2616_/A sky130_fd_sc_hd__and2_1
X_1428_ _1428_/A vssd1 vssd1 vccd1 vccd1 _1440_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2477_ _2481_/A vssd1 vssd1 vccd1 vccd1 _2477_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2546_ _2546_/A _2546_/B vssd1 vssd1 vccd1 vccd1 _2547_/A sky130_fd_sc_hd__and2_1
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1359_ _2751_/Q _2750_/Q _1359_/C _1359_/D vssd1 vssd1 vccd1 vccd1 _1360_/B sky130_fd_sc_hd__or4_4
XFILLER_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2400_ _2709_/Q _2710_/Q _2400_/C vssd1 vssd1 vccd1 vccd1 _2404_/B sky130_fd_sc_hd__and3_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2262_ _2262_/A vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__clkinv_2
X_2331_ _2685_/Q _2332_/C _2686_/Q vssd1 vssd1 vccd1 vccd1 _2333_/A sky130_fd_sc_hd__a21oi_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2193_ input1/X vssd1 vssd1 vccd1 vccd1 _2571_/A sky130_fd_sc_hd__inv_2
X_1977_ _1978_/A _1977_/B vssd1 vssd1 vccd1 vccd1 _1977_/Y sky130_fd_sc_hd__xnor2_1
X_2529_ _2788_/Q vssd1 vssd1 vccd1 vccd1 _2590_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1900_ _1900_/A _1900_/B vssd1 vssd1 vccd1 vccd1 _1901_/C sky130_fd_sc_hd__nor2_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1831_ _2052_/B vssd1 vssd1 vccd1 vccd1 _1831_/Y sky130_fd_sc_hd__clkinv_2
X_1693_ _1902_/B _1713_/C vssd1 vssd1 vccd1 vccd1 _1719_/A sky130_fd_sc_hd__xor2_2
X_1762_ _1762_/A vssd1 vssd1 vccd1 vccd1 _1792_/A sky130_fd_sc_hd__clkbuf_2
X_2314_ _2678_/Q _2314_/B vssd1 vssd1 vccd1 vccd1 _2318_/C sky130_fd_sc_hd__and2_1
X_2245_ _2245_/A vssd1 vssd1 vccd1 vccd1 _2773_/D sky130_fd_sc_hd__clkbuf_1
X_2176_ _2773_/Q vssd1 vssd1 vccd1 vccd1 _2527_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2030_ _2030_/A _2034_/A vssd1 vssd1 vccd1 vccd1 _2031_/B sky130_fd_sc_hd__or2_1
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1745_ _1745_/A _1745_/B vssd1 vssd1 vccd1 vccd1 _1793_/A sky130_fd_sc_hd__xor2_2
X_2794_ _2805_/CLK _2794_/D vssd1 vssd1 vccd1 vccd1 _2794_/Q sky130_fd_sc_hd__dfxtp_1
X_1814_ _1842_/B vssd1 vssd1 vccd1 vccd1 _1917_/A sky130_fd_sc_hd__clkbuf_2
X_1676_ _1901_/B _1679_/B vssd1 vssd1 vccd1 vccd1 _1685_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2228_ _2228_/A _2233_/B vssd1 vssd1 vccd1 vccd1 _2229_/A sky130_fd_sc_hd__or2b_2
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2159_ _2159_/A vssd1 vssd1 vccd1 vccd1 _2159_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1392_ _1392_/A _1555_/A vssd1 vssd1 vccd1 vccd1 _1403_/A sky130_fd_sc_hd__xnor2_2
X_1461_ _1461_/A vssd1 vssd1 vccd1 vccd1 _1470_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1530_ _1530_/A _1544_/A vssd1 vssd1 vccd1 vccd1 _1539_/B sky130_fd_sc_hd__xor2_2
X_2013_ _2013_/A _2013_/B vssd1 vssd1 vccd1 vccd1 _2013_/Y sky130_fd_sc_hd__xnor2_1
X_1728_ _1728_/A _1728_/B vssd1 vssd1 vccd1 vccd1 _1728_/X sky130_fd_sc_hd__or2_1
X_2777_ _2788_/CLK _2777_/D vssd1 vssd1 vccd1 vccd1 _2777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ _1650_/Y _1665_/A _1656_/Y _1658_/X vssd1 vssd1 vccd1 vccd1 _1661_/C sky130_fd_sc_hd__o31ai_4
XFILLER_37_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2700_ _2806_/CLK _2700_/D vssd1 vssd1 vccd1 vccd1 _2700_/Q sky130_fd_sc_hd__dfxtp_1
X_2562_ _2562_/A vssd1 vssd1 vccd1 vccd1 _2794_/D sky130_fd_sc_hd__clkbuf_1
X_2631_ _2803_/Q _2617_/X _2630_/X _2358_/X vssd1 vssd1 vccd1 vccd1 _2803_/D sky130_fd_sc_hd__o211a_1
X_1444_ _1444_/A _1444_/B _1571_/B vssd1 vssd1 vccd1 vccd1 _1456_/B sky130_fd_sc_hd__and3_1
X_1375_ _1375_/A _1410_/B _1375_/C vssd1 vssd1 vccd1 vccd1 _1549_/B sky130_fd_sc_hd__or3_1
X_1513_ _1749_/A _2057_/A _1522_/B vssd1 vssd1 vccd1 vccd1 _1514_/B sky130_fd_sc_hd__a21boi_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2493_ _2494_/A vssd1 vssd1 vccd1 vccd1 _2493_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _1983_/X _1991_/Y _1993_/S vssd1 vssd1 vccd1 vccd1 _2029_/B sky130_fd_sc_hd__mux2_1
X_2614_ _2800_/Q _2597_/X _2613_/X _2601_/A vssd1 vssd1 vccd1 vccd1 _2615_/B sky130_fd_sc_hd__a22o_1
X_2545_ _2791_/Q _2544_/X _2550_/S vssd1 vssd1 vccd1 vccd1 _2546_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1427_ _1428_/A _1433_/A _1433_/B _1430_/A _1430_/B vssd1 vssd1 vccd1 vccd1 _1557_/C
+ sky130_fd_sc_hd__o311ai_4
X_1358_ _2749_/Q _2748_/Q vssd1 vssd1 vccd1 vccd1 _1359_/D sky130_fd_sc_hd__or2_1
X_2476_ _2489_/A vssd1 vssd1 vccd1 vccd1 _2481_/A sky130_fd_sc_hd__buf_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2330_ _2685_/Q _2332_/C vssd1 vssd1 vccd1 vccd1 _2685_/D sky130_fd_sc_hd__xor2_1
X_2261_ _2663_/Q _2262_/A vssd1 vssd1 vccd1 vccd1 _2273_/B sky130_fd_sc_hd__or2_1
X_2192_ _2192_/A vssd1 vssd1 vccd1 vccd1 _2772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1976_ _1976_/A vssd1 vssd1 vccd1 vccd1 _1978_/A sky130_fd_sc_hd__inv_2
X_2528_ _2525_/Y _2527_/Y _2511_/A vssd1 vssd1 vccd1 vccd1 _2787_/D sky130_fd_sc_hd__a21oi_1
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2459_ _2463_/A vssd1 vssd1 vccd1 vccd1 _2459_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2823__26 vssd1 vssd1 vccd1 vccd1 _2823__26/HI o_io_oeb[12] sky130_fd_sc_hd__conb_1
XFILLER_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1830_ _1887_/A vssd1 vssd1 vccd1 vccd1 _2041_/A sky130_fd_sc_hd__clkbuf_2
X_1761_ _1903_/B _1775_/A vssd1 vssd1 vccd1 vccd1 _1793_/C sky130_fd_sc_hd__or2_1
X_2313_ _2678_/Q _2314_/B vssd1 vssd1 vccd1 vccd1 _2315_/A sky130_fd_sc_hd__nor2_1
X_1692_ _1714_/A _1704_/A _1704_/B _1739_/A _1691_/Y vssd1 vssd1 vccd1 vccd1 _1713_/C
+ sky130_fd_sc_hd__o41a_2
X_2175_ _2445_/A vssd1 vssd1 vccd1 vccd1 _2511_/A sky130_fd_sc_hd__clkbuf_2
X_2244_ _2244_/A _2636_/A vssd1 vssd1 vccd1 vccd1 _2245_/A sky130_fd_sc_hd__and2_1
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ _1976_/A _1978_/B vssd1 vssd1 vccd1 vccd1 _1971_/A sky130_fd_sc_hd__or2_1
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1744_ _1744_/A _1758_/A _1760_/B vssd1 vssd1 vccd1 vccd1 _1745_/B sky130_fd_sc_hd__and3_1
XFILLER_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2793_ _2793_/CLK _2793_/D vssd1 vssd1 vccd1 vccd1 _2793_/Q sky130_fd_sc_hd__dfxtp_1
X_1813_ _1808_/X _1810_/X _1812_/X vssd1 vssd1 vccd1 vccd1 _1842_/B sky130_fd_sc_hd__o21ai_2
X_1675_ _1675_/A vssd1 vssd1 vccd1 vccd1 _1714_/A sky130_fd_sc_hd__inv_2
X_2089_ _2089_/A vssd1 vssd1 vccd1 vccd1 _2089_/Y sky130_fd_sc_hd__inv_2
X_2227_ _2227_/A _2227_/B _2227_/C vssd1 vssd1 vccd1 vccd1 _2233_/B sky130_fd_sc_hd__or3_2
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2158_ _2137_/X _2156_/Y _2157_/X _2146_/X _2157_/A vssd1 vssd1 vccd1 vccd1 _2732_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1460_ _1470_/B vssd1 vssd1 vccd1 vccd1 _1590_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1391_ _1391_/A _1391_/B vssd1 vssd1 vccd1 vccd1 _1391_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2012_ _2170_/A _2767_/Q _2010_/Y _2011_/X vssd1 vssd1 vccd1 vccd1 _2767_/D sky130_fd_sc_hd__o22a_1
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1658_ _1658_/A _1658_/B vssd1 vssd1 vccd1 vccd1 _1658_/X sky130_fd_sc_hd__xor2_2
X_1727_ _1722_/A _1720_/B _1696_/A vssd1 vssd1 vccd1 vccd1 _1728_/B sky130_fd_sc_hd__a21oi_1
X_2776_ _2783_/CLK _2776_/D vssd1 vssd1 vccd1 vccd1 _2776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1589_ _1619_/C _1586_/X _1587_/Y _1588_/Y vssd1 vssd1 vccd1 vccd1 _1589_/X sky130_fd_sc_hd__a211o_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1512_ _1512_/A _1512_/B vssd1 vssd1 vccd1 vccd1 _1522_/B sky130_fd_sc_hd__nand2_1
X_2561_ _2569_/A _2561_/B vssd1 vssd1 vccd1 vccd1 _2562_/A sky130_fd_sc_hd__and2_1
X_2492_ _2494_/A vssd1 vssd1 vccd1 vccd1 _2492_/Y sky130_fd_sc_hd__inv_2
X_2630_ _2802_/Q _2249_/A _2629_/X _2244_/A _2625_/X vssd1 vssd1 vccd1 vccd1 _2630_/X
+ sky130_fd_sc_hd__a221o_1
X_1443_ _1571_/A _1571_/B _1444_/A vssd1 vssd1 vccd1 vccd1 _1456_/A sky130_fd_sc_hd__a21oi_1
X_1374_ _2758_/Q _1374_/B _1374_/C vssd1 vssd1 vccd1 vccd1 _1375_/C sky130_fd_sc_hd__or3_1
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2759_ _2759_/CLK _2759_/D _2481_/Y vssd1 vssd1 vccd1 vccd1 _2759_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1992_ _1992_/A _1992_/B vssd1 vssd1 vccd1 vccd1 _1993_/S sky130_fd_sc_hd__nand2_1
X_2475_ _2475_/A vssd1 vssd1 vccd1 vccd1 _2475_/Y sky130_fd_sc_hd__inv_2
X_2613_ _2799_/Q _2598_/X _2612_/X vssd1 vssd1 vccd1 vccd1 _2613_/X sky130_fd_sc_hd__a21bo_1
X_2544_ _2763_/Q _2790_/Q _2553_/S vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1426_ _1551_/A _1551_/B _1409_/Y _1424_/A vssd1 vssd1 vccd1 vccd1 _1430_/B sky130_fd_sc_hd__a211o_1
X_1357_ _1458_/A vssd1 vssd1 vccd1 vccd1 _1474_/A sky130_fd_sc_hd__inv_2
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2260_ _2663_/Q _2262_/A vssd1 vssd1 vccd1 vccd1 _2275_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2191_ _2489_/A _2776_/Q _2190_/X vssd1 vssd1 vccd1 vccd1 _2192_/A sky130_fd_sc_hd__or3b_1
XFILLER_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _1975_/A vssd1 vssd1 vccd1 vccd1 _1975_/Y sky130_fd_sc_hd__inv_2
X_1409_ _1409_/A _1579_/B vssd1 vssd1 vccd1 vccd1 _1409_/Y sky130_fd_sc_hd__xnor2_2
X_2458_ _2470_/A vssd1 vssd1 vccd1 vccd1 _2463_/A sky130_fd_sc_hd__buf_2
X_2527_ _2527_/A _2632_/B vssd1 vssd1 vccd1 vccd1 _2527_/Y sky130_fd_sc_hd__nand2_1
X_2389_ _2705_/Q _2390_/B vssd1 vssd1 vccd1 vccd1 _2393_/C sky130_fd_sc_hd__and2_1
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1691_ _1691_/A _1691_/B vssd1 vssd1 vccd1 vccd1 _1691_/Y sky130_fd_sc_hd__xnor2_1
X_1760_ _1903_/A _1760_/B vssd1 vssd1 vccd1 vccd1 _1775_/A sky130_fd_sc_hd__xor2_4
X_2312_ _2312_/A _2314_/B vssd1 vssd1 vccd1 vccd1 _2677_/D sky130_fd_sc_hd__nor2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2174_ input1/X vssd1 vssd1 vccd1 vccd1 _2445_/A sky130_fd_sc_hd__clkbuf_2
X_2243_ _2571_/A vssd1 vssd1 vccd1 vccd1 _2636_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1958_ _1963_/A _1960_/C vssd1 vssd1 vccd1 vccd1 _1978_/B sky130_fd_sc_hd__xor2_1
X_1889_ _1890_/B _1889_/B _1888_/X vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__or3b_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1674_ _1674_/A _1674_/B vssd1 vssd1 vccd1 vccd1 _1675_/A sky130_fd_sc_hd__nor2_1
X_1743_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1744_/A sky130_fd_sc_hd__clkbuf_2
X_2792_ _2793_/CLK _2792_/D vssd1 vssd1 vccd1 vccd1 _2792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1812_ _1811_/A _1811_/Y _1812_/S vssd1 vssd1 vccd1 vccd1 _1812_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2226_ _2226_/A vssd1 vssd1 vccd1 vccd1 _2226_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2088_ _2113_/A vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__clkbuf_2
X_2157_ _2157_/A _2159_/A vssd1 vssd1 vccd1 vccd1 _2157_/X sky130_fd_sc_hd__or2_1
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1390_ _1390_/A _1394_/B _1549_/A vssd1 vssd1 vccd1 vccd1 _1391_/B sky130_fd_sc_hd__or3b_1
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2011_ _1915_/B _1923_/X _1996_/Y _2003_/A vssd1 vssd1 vccd1 vccd1 _2011_/X sky130_fd_sc_hd__a31o_1
X_1588_ _1620_/A vssd1 vssd1 vccd1 vccd1 _1588_/Y sky130_fd_sc_hd__inv_2
X_1657_ _1639_/D _1642_/B _1645_/Y _1655_/A vssd1 vssd1 vccd1 vccd1 _1658_/B sky130_fd_sc_hd__a22o_1
X_1726_ _1721_/S _1720_/B _1696_/A _1722_/A vssd1 vssd1 vccd1 vccd1 _1728_/A sky130_fd_sc_hd__o211a_1
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2775_ _2809_/CLK _2775_/D vssd1 vssd1 vccd1 vccd1 _2775_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _2657_/Q _2234_/B vssd1 vssd1 vccd1 vccd1 _2235_/B sky130_fd_sc_hd__nor2_4
XFILLER_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1442_ _1431_/C _1563_/B _1441_/X vssd1 vssd1 vccd1 vccd1 _1571_/B sky130_fd_sc_hd__o21a_1
X_1511_ _2741_/Q _2740_/Q _1805_/B _1511_/D vssd1 vssd1 vccd1 vccd1 _1512_/B sky130_fd_sc_hd__or4_1
X_2560_ _2794_/Q _2559_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2561_/B sky130_fd_sc_hd__mux2_1
X_2491_ _2494_/A vssd1 vssd1 vccd1 vccd1 _2491_/Y sky130_fd_sc_hd__inv_2
X_1373_ _1373_/A vssd1 vssd1 vccd1 vccd1 _1375_/A sky130_fd_sc_hd__clkinv_2
X_2758_ _2758_/CLK _2758_/D _2480_/Y vssd1 vssd1 vccd1 vccd1 _2758_/Q sky130_fd_sc_hd__dfrtp_1
X_2689_ _2760_/CLK _2689_/D vssd1 vssd1 vccd1 vccd1 _2689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1709_ _1902_/B _1713_/C vssd1 vssd1 vccd1 vccd1 _1710_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1991_ _1991_/A _1991_/B vssd1 vssd1 vccd1 vccd1 _1991_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2612_ _2622_/A _2633_/A _2622_/C _2576_/A vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__or4b_1
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1425_ _1424_/A _1551_/B _1409_/Y vssd1 vssd1 vccd1 vccd1 _1430_/A sky130_fd_sc_hd__o21ai_2
X_2474_ _2475_/A vssd1 vssd1 vccd1 vccd1 _2474_/Y sky130_fd_sc_hd__inv_2
X_2543_ _2543_/A vssd1 vssd1 vccd1 vccd1 _2790_/D sky130_fd_sc_hd__clkbuf_1
X_1356_ _2749_/Q _1356_/B vssd1 vssd1 vccd1 vccd1 _1458_/A sky130_fd_sc_hd__xnor2_2
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2190_ _2771_/Q _2772_/Q vssd1 vssd1 vccd1 vccd1 _2190_/X sky130_fd_sc_hd__or2b_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1974_ _1991_/B _1974_/B vssd1 vssd1 vccd1 vccd1 _1992_/A sky130_fd_sc_hd__and2_1
X_1408_ _1412_/B _1413_/S _1412_/A vssd1 vssd1 vccd1 vccd1 _1579_/B sky130_fd_sc_hd__a21o_2
X_2388_ _2390_/B _2388_/B vssd1 vssd1 vccd1 vccd1 _2704_/D sky130_fd_sc_hd__nor2_1
X_2457_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2457_/Y sky130_fd_sc_hd__inv_2
X_2526_ _2787_/Q _2581_/B vssd1 vssd1 vccd1 vccd1 _2632_/B sky130_fd_sc_hd__nor2_2
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1339_ _1510_/A _1829_/B _1339_/C _1511_/D vssd1 vssd1 vccd1 vccd1 _1360_/A sky130_fd_sc_hd__or4_2
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2814__17 vssd1 vssd1 vccd1 vccd1 _2814__17/HI o_io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1690_ _1688_/A _1711_/A _1675_/A _1688_/B _1674_/A vssd1 vssd1 vccd1 vccd1 _1691_/B
+ sky130_fd_sc_hd__a41o_1
X_2311_ _2676_/Q _2677_/Q _2311_/C vssd1 vssd1 vccd1 vccd1 _2314_/B sky130_fd_sc_hd__and3_1
X_2242_ _2242_/A vssd1 vssd1 vccd1 vccd1 _2244_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2173_ _2208_/A vssd1 vssd1 vccd1 vccd1 _2657_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ _1960_/C vssd1 vssd1 vccd1 vccd1 _2022_/A sky130_fd_sc_hd__buf_2
X_1888_ _2163_/A _1888_/B vssd1 vssd1 vccd1 vccd1 _1888_/X sky130_fd_sc_hd__xor2_1
X_2509_ _2781_/Q _2510_/C _2782_/Q vssd1 vssd1 vccd1 vccd1 _2511_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2791_ _2793_/CLK _2791_/D vssd1 vssd1 vccd1 vccd1 _2791_/Q sky130_fd_sc_hd__dfxtp_1
X_1811_ _1811_/A _1904_/A vssd1 vssd1 vccd1 vccd1 _1811_/Y sky130_fd_sc_hd__nand2_1
X_1673_ _1672_/X _1679_/B _1662_/Y _1661_/X vssd1 vssd1 vccd1 vccd1 _1674_/B sky130_fd_sc_hd__a211oi_1
XFILLER_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1742_ _1767_/B _1742_/B vssd1 vssd1 vccd1 vccd1 _1793_/B sky130_fd_sc_hd__xnor2_1
X_2225_ _2221_/A _2225_/B _2225_/C vssd1 vssd1 vccd1 vccd1 _2226_/A sky130_fd_sc_hd__and3b_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2087_ _2083_/B _2085_/Y _2065_/A _2086_/X vssd1 vssd1 vccd1 vccd1 _2755_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2156_ _2157_/A _2159_/A vssd1 vssd1 vccd1 vccd1 _2156_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2010_ _1923_/X _1996_/Y _1915_/B vssd1 vssd1 vccd1 vccd1 _2010_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1725_ _2739_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1756_/B sky130_fd_sc_hd__xnor2_1
X_2774_ _2783_/CLK _2774_/D vssd1 vssd1 vccd1 vccd1 _2774_/Q sky130_fd_sc_hd__dfxtp_1
X_1587_ _1619_/A _1587_/B vssd1 vssd1 vccd1 vccd1 _1587_/Y sky130_fd_sc_hd__nor2_1
X_1656_ _1669_/A _1682_/A vssd1 vssd1 vccd1 vccd1 _1656_/Y sky130_fd_sc_hd__nand2_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _2208_/A _2658_/Q vssd1 vssd1 vccd1 vccd1 _2235_/A sky130_fd_sc_hd__nor2_2
XFILLER_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2139_ _2142_/A _2144_/A _2055_/A vssd1 vssd1 vccd1 vccd1 _2139_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1441_ _1440_/Y _1409_/Y _1433_/Y _1557_/B vssd1 vssd1 vccd1 vccd1 _1441_/X sky130_fd_sc_hd__a31o_1
X_1510_ _1510_/A _1829_/B vssd1 vssd1 vccd1 vccd1 _1805_/B sky130_fd_sc_hd__or2_2
XFILLER_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2490_ _2494_/A vssd1 vssd1 vccd1 vccd1 _2490_/Y sky130_fd_sc_hd__inv_2
X_1372_ _1365_/Y _1367_/Y _1390_/A vssd1 vssd1 vccd1 vccd1 _1549_/A sky130_fd_sc_hd__a21o_1
X_2688_ _2727_/CLK _2688_/D vssd1 vssd1 vccd1 vccd1 _2688_/Q sky130_fd_sc_hd__dfxtp_1
X_2757_ _2757_/CLK _2757_/D _2479_/Y vssd1 vssd1 vccd1 vccd1 _2757_/Q sky130_fd_sc_hd__dfrtp_1
X_1708_ _1719_/A _1731_/A vssd1 vssd1 vccd1 vccd1 _1734_/A sky130_fd_sc_hd__nand2_1
X_1639_ _1644_/A _1644_/B _1642_/B _1639_/D vssd1 vssd1 vccd1 vccd1 _1639_/X sky130_fd_sc_hd__and4bb_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1990_ _1985_/X _1987_/Y _1988_/X _1989_/Y _1992_/A vssd1 vssd1 vccd1 vccd1 _2029_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_13_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2542_ _2546_/A _2542_/B vssd1 vssd1 vccd1 vccd1 _2543_/A sky130_fd_sc_hd__and2_1
X_2611_ _2611_/A _2611_/B vssd1 vssd1 vccd1 vccd1 _2633_/A sky130_fd_sc_hd__or2_1
X_1424_ _1424_/A _1551_/A _1551_/B vssd1 vssd1 vccd1 vccd1 _1433_/B sky130_fd_sc_hd__and3_1
X_1355_ _1334_/A _2748_/Q _1454_/B vssd1 vssd1 vccd1 vccd1 _1356_/B sky130_fd_sc_hd__a21o_1
X_2473_ _2475_/A vssd1 vssd1 vccd1 vccd1 _2473_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2809_ _2809_/CLK _2809_/D vssd1 vssd1 vccd1 vccd1 _2809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ _1971_/A _1977_/B _1971_/B vssd1 vssd1 vccd1 vccd1 _1974_/B sky130_fd_sc_hd__a21o_1
X_2525_ _2525_/A _2525_/B vssd1 vssd1 vccd1 vccd1 _2525_/Y sky130_fd_sc_hd__nand2_1
X_1407_ _1409_/A _1407_/B _1407_/C vssd1 vssd1 vccd1 vccd1 _1412_/B sky130_fd_sc_hd__or3_1
X_2387_ _2703_/Q _2386_/C _2704_/Q vssd1 vssd1 vccd1 vccd1 _2388_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2456_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2456_/Y sky130_fd_sc_hd__inv_2
X_1338_ _2739_/Q _2738_/Q _2737_/Q _2736_/Q vssd1 vssd1 vccd1 vccd1 _1511_/D sky130_fd_sc_hd__or4_1
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2310_ _2676_/Q _2311_/C _2677_/Q vssd1 vssd1 vccd1 vccd1 _2312_/A sky130_fd_sc_hd__a21oi_1
X_2172_ _2657_/Q vssd1 vssd1 vccd1 vccd1 _2208_/A sky130_fd_sc_hd__inv_2
X_2241_ _2576_/A vssd1 vssd1 vccd1 vccd1 _2242_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1887_ _1887_/A _1887_/B vssd1 vssd1 vccd1 vccd1 _1888_/B sky130_fd_sc_hd__nand2_1
X_1956_ _1943_/X _1983_/A _1965_/B _1965_/C _1955_/X vssd1 vssd1 vccd1 vccd1 _1960_/C
+ sky130_fd_sc_hd__a41o_1
X_2508_ _2508_/A vssd1 vssd1 vccd1 vccd1 _2781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2439_ _2726_/Q _2439_/B vssd1 vssd1 vccd1 vccd1 _2440_/B sky130_fd_sc_hd__or2_1
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2790_ _2793_/CLK _2790_/D vssd1 vssd1 vccd1 vccd1 _2790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1810_ _1811_/A _1784_/X _1809_/X vssd1 vssd1 vccd1 vccd1 _1810_/X sky130_fd_sc_hd__o21a_1
X_1741_ _1767_/C _1760_/B vssd1 vssd1 vccd1 vccd1 _1742_/B sky130_fd_sc_hd__nand2_1
X_1672_ _1672_/A _1680_/A vssd1 vssd1 vccd1 vccd1 _1672_/X sky130_fd_sc_hd__or2_1
XFILLER_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2224_ _2227_/A _2227_/B vssd1 vssd1 vccd1 vccd1 _2225_/C sky130_fd_sc_hd__and2b_1
X_2155_ _2052_/A _2070_/X _2073_/X _2154_/Y vssd1 vssd1 vccd1 vccd1 _2733_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2086_ _2099_/A vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1939_ _1946_/B vssd1 vssd1 vccd1 vccd1 _2018_/A sky130_fd_sc_hd__buf_2
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_14_0_i_clk clkbuf_3_7_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _2760_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1724_ _2738_/Q _2055_/B _2736_/Q _1805_/B _1749_/A vssd1 vssd1 vccd1 vccd1 _1725_/B
+ sky130_fd_sc_hd__o41a_1
X_2773_ _2788_/CLK _2773_/D vssd1 vssd1 vccd1 vccd1 _2773_/Q sky130_fd_sc_hd__dfxtp_1
X_1586_ _1573_/A _1619_/A _1619_/B vssd1 vssd1 vccd1 vccd1 _1586_/X sky130_fd_sc_hd__mux2_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ _1655_/A _1655_/B vssd1 vssd1 vccd1 vccd1 _1682_/A sky130_fd_sc_hd__nor2_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _2227_/A _2227_/B vssd1 vssd1 vccd1 vccd1 _2222_/A sky130_fd_sc_hd__nor2_1
X_2138_ _2138_/A vssd1 vssd1 vccd1 vccd1 _2138_/Y sky130_fd_sc_hd__inv_2
X_2069_ _2068_/A _1327_/B _2692_/D _2170_/B vssd1 vssd1 vccd1 vccd1 _2146_/A sky130_fd_sc_hd__a211o_1
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1440_ _1440_/A vssd1 vssd1 vccd1 vccd1 _1440_/Y sky130_fd_sc_hd__inv_2
X_1371_ _2075_/A _1371_/B vssd1 vssd1 vccd1 vccd1 _1390_/A sky130_fd_sc_hd__xnor2_1
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2687_ _2727_/CLK _2687_/D vssd1 vssd1 vccd1 vccd1 _2687_/Q sky130_fd_sc_hd__dfxtp_1
X_1638_ _1638_/A _1638_/B vssd1 vssd1 vccd1 vccd1 _1639_/D sky130_fd_sc_hd__nor2_1
X_1707_ _1737_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1733_/A sky130_fd_sc_hd__and2_1
X_2756_ _2802_/CLK _2756_/D _2478_/Y vssd1 vssd1 vccd1 vccd1 _2756_/Q sky130_fd_sc_hd__dfrtp_2
X_1569_ _1576_/A _1569_/B vssd1 vssd1 vccd1 vccd1 _1620_/A sky130_fd_sc_hd__xnor2_2
XFILLER_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2472_ _2475_/A vssd1 vssd1 vccd1 vccd1 _2472_/Y sky130_fd_sc_hd__inv_2
X_2541_ _2790_/Q _2540_/X _2550_/S vssd1 vssd1 vccd1 vccd1 _2542_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2610_ _2610_/A _2610_/B vssd1 vssd1 vccd1 vccd1 _2611_/B sky130_fd_sc_hd__and2_1
X_1423_ _1551_/A _1551_/B _1424_/A vssd1 vssd1 vccd1 vccd1 _1433_/A sky130_fd_sc_hd__a21oi_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1354_ _1341_/B _1359_/C _1410_/A vssd1 vssd1 vccd1 vccd1 _1454_/B sky130_fd_sc_hd__o21a_1
XFILLER_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2808_ _2809_/CLK _2808_/D vssd1 vssd1 vccd1 vccd1 _2808_/Q sky130_fd_sc_hd__dfxtp_1
X_2739_ _2759_/CLK _2739_/D _2457_/Y vssd1 vssd1 vccd1 vccd1 _2739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _1972_/A _1978_/C vssd1 vssd1 vccd1 vccd1 _1991_/B sky130_fd_sc_hd__nand2_1
X_2455_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2455_/Y sky130_fd_sc_hd__inv_2
X_2524_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2525_/A sky130_fd_sc_hd__clkbuf_2
X_1406_ _1406_/A vssd1 vssd1 vccd1 vccd1 _1409_/A sky130_fd_sc_hd__inv_2
X_2386_ _2703_/Q _2704_/Q _2386_/C vssd1 vssd1 vccd1 vccd1 _2390_/B sky130_fd_sc_hd__and3_1
X_1337_ _2743_/Q _2742_/Q _2741_/Q _2740_/Q vssd1 vssd1 vccd1 vccd1 _1339_/C sky130_fd_sc_hd__or4_1
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2171_ _2171_/A vssd1 vssd1 vccd1 vccd1 _2695_/D sky130_fd_sc_hd__clkbuf_1
X_2240_ _2777_/Q vssd1 vssd1 vccd1 vccd1 _2576_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1955_ _1936_/B _1948_/Y _1951_/Y _1954_/Y vssd1 vssd1 vccd1 vccd1 _1955_/X sky130_fd_sc_hd__o31a_1
X_1886_ _2730_/Q vssd1 vssd1 vccd1 vccd1 _2163_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2438_ _2726_/Q _2439_/B vssd1 vssd1 vccd1 vccd1 _2442_/B sky130_fd_sc_hd__nand2_1
X_2507_ _2636_/A _2507_/B _2507_/C _2507_/D vssd1 vssd1 vccd1 vccd1 _2508_/A sky130_fd_sc_hd__and4_1
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2369_ _2697_/Q _2696_/Q _2698_/Q vssd1 vssd1 vccd1 vccd1 _2373_/C sky130_fd_sc_hd__and3_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_10_0_i_clk clkbuf_3_5_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _2726_/CLK sky130_fd_sc_hd__clkbuf_2
X_1671_ _1671_/A _1679_/B vssd1 vssd1 vccd1 vccd1 _1674_/A sky130_fd_sc_hd__and2_1
X_1740_ _1767_/A _1767_/B _1767_/C _1762_/A _1763_/D vssd1 vssd1 vccd1 vccd1 _1760_/B
+ sky130_fd_sc_hd__a41o_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2085_ _2065_/A _2089_/A _2043_/X vssd1 vssd1 vccd1 vccd1 _2085_/Y sky130_fd_sc_hd__o21ai_1
X_2223_ _2223_/A vssd1 vssd1 vccd1 vccd1 _2223_/X sky130_fd_sc_hd__clkbuf_1
X_2154_ _2154_/A _2154_/B vssd1 vssd1 vccd1 vccd1 _2154_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1938_ _1925_/Y _1941_/A _1951_/A _1951_/B _1937_/X vssd1 vssd1 vccd1 vccd1 _1946_/B
+ sky130_fd_sc_hd__a41oi_2
X_1869_ _1870_/A _1869_/B vssd1 vssd1 vccd1 vccd1 _1869_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1654_ _1636_/A _1640_/X _1643_/Y vssd1 vssd1 vccd1 vccd1 _1655_/B sky130_fd_sc_hd__a21oi_1
X_1723_ _2737_/Q vssd1 vssd1 vccd1 vccd1 _2055_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2772_ _2783_/CLK _2772_/D vssd1 vssd1 vccd1 vccd1 _2772_/Q sky130_fd_sc_hd__dfxtp_1
X_1585_ _1585_/A vssd1 vssd1 vccd1 vccd1 _1619_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2808_/Q _2234_/B _2205_/X vssd1 vssd1 vccd1 vccd1 _2227_/B sky130_fd_sc_hd__o21ai_2
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2068_ _2068_/A _2068_/B vssd1 vssd1 vccd1 vccd1 _2170_/B sky130_fd_sc_hd__nor2_1
X_2137_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1370_ _1360_/A _1360_/B _1374_/B _1374_/C _1373_/A vssd1 vssd1 vccd1 vccd1 _1371_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1637_ _1637_/A _1644_/A vssd1 vssd1 vccd1 vccd1 _1637_/Y sky130_fd_sc_hd__xnor2_1
X_2686_ _2727_/CLK _2686_/D vssd1 vssd1 vccd1 vccd1 _2686_/Q sky130_fd_sc_hd__dfxtp_1
X_2755_ _2757_/CLK _2755_/D _2477_/Y vssd1 vssd1 vccd1 vccd1 _2755_/Q sky130_fd_sc_hd__dfrtp_1
X_1706_ _1704_/B _1691_/Y _1704_/A vssd1 vssd1 vccd1 vccd1 _1707_/B sky130_fd_sc_hd__o21ai_1
X_1568_ _1581_/B _1577_/C vssd1 vssd1 vccd1 vccd1 _1569_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1499_ _1499_/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1499_/Y sky130_fd_sc_hd__nand2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2471_ _2475_/A vssd1 vssd1 vccd1 vccd1 _2471_/Y sky130_fd_sc_hd__inv_2
X_1422_ _2063_/A _1422_/B vssd1 vssd1 vccd1 vccd1 _1424_/A sky130_fd_sc_hd__xnor2_2
X_2540_ _2762_/Q _2789_/Q _2553_/S vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1353_ _2747_/Q _2746_/Q _2745_/Q _2744_/Q vssd1 vssd1 vccd1 vccd1 _1359_/C sky130_fd_sc_hd__or4_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2738_ _2759_/CLK _2738_/D _2456_/Y vssd1 vssd1 vccd1 vccd1 _2738_/Q sky130_fd_sc_hd__dfrtp_1
X_2807_ _2807_/CLK _2807_/D vssd1 vssd1 vccd1 vccd1 _2807_/Q sky130_fd_sc_hd__dfxtp_1
X_2669_ _2727_/CLK _2669_/D vssd1 vssd1 vccd1 vccd1 _2669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1971_ _1971_/A _1971_/B vssd1 vssd1 vccd1 vccd1 _1972_/A sky130_fd_sc_hd__and2_1
X_1405_ _1405_/A _1405_/B vssd1 vssd1 vccd1 vccd1 _1405_/X sky130_fd_sc_hd__or2_1
X_2385_ _2703_/Q _2386_/C vssd1 vssd1 vccd1 vccd1 _2703_/D sky130_fd_sc_hd__xor2_1
X_2454_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2454_/Y sky130_fd_sc_hd__inv_2
X_2523_ _2527_/A _2521_/X _2546_/A _2525_/B vssd1 vssd1 vccd1 vccd1 _2786_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1336_ _2731_/Q _2730_/Q _2729_/Q _2728_/Q vssd1 vssd1 vccd1 vccd1 _1829_/B sky130_fd_sc_hd__or4_4
Xinput1 i_reset vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2170_ _2170_/A _2170_/B vssd1 vssd1 vccd1 vccd1 _2171_/A sky130_fd_sc_hd__or2_1
X_1954_ _1948_/Y _1951_/Y _2018_/A _1953_/Y vssd1 vssd1 vccd1 vccd1 _1954_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1885_ _1875_/A _1985_/A vssd1 vssd1 vccd1 vccd1 _1889_/B sky130_fd_sc_hd__and2b_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2437_ _2439_/B _2437_/B vssd1 vssd1 vccd1 vccd1 _2725_/D sky130_fd_sc_hd__nor2_1
X_2368_ _2697_/Q _2696_/Q _2698_/Q vssd1 vssd1 vccd1 vccd1 _2370_/A sky130_fd_sc_hd__a21oi_1
X_2506_ _2781_/Q _2510_/C vssd1 vssd1 vccd1 vccd1 _2507_/D sky130_fd_sc_hd__nand2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2299_ _2672_/Q _2671_/Q _2299_/C vssd1 vssd1 vccd1 vccd1 _2307_/D sky130_fd_sc_hd__and3_1
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1670_ _1682_/A _1671_/A _1691_/A _1669_/X vssd1 vssd1 vccd1 vccd1 _1679_/B sky130_fd_sc_hd__a31o_1
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2222_ _2222_/A _2222_/B _2227_/C vssd1 vssd1 vccd1 vccd1 _2223_/A sky130_fd_sc_hd__and3_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ _2073_/X _2082_/Y _2083_/X _2077_/X _2083_/A vssd1 vssd1 vccd1 vccd1 _2756_/D
+ sky130_fd_sc_hd__a32o_1
X_2153_ _2157_/A _2159_/A _2052_/A vssd1 vssd1 vccd1 vccd1 _2154_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1937_ _1934_/X _1953_/A _1936_/X _1935_/B vssd1 vssd1 vccd1 vccd1 _1937_/X sky130_fd_sc_hd__o2bb2a_1
X_1868_ _1870_/B _1963_/A vssd1 vssd1 vccd1 vccd1 _1869_/B sky130_fd_sc_hd__nand2_1
X_1799_ _1910_/A _1910_/B vssd1 vssd1 vccd1 vccd1 _1803_/A sky130_fd_sc_hd__xor2_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2771_ _2809_/CLK _2771_/D _2495_/Y vssd1 vssd1 vccd1 vccd1 _2771_/Q sky130_fd_sc_hd__dfrtp_1
X_1584_ _1591_/B vssd1 vssd1 vccd1 vccd1 _1619_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_1653_ _1647_/X _1640_/X _1643_/Y _1636_/A vssd1 vssd1 vccd1 vccd1 _1655_/A sky130_fd_sc_hd__o211a_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _1722_/A _1731_/A vssd1 vssd1 vccd1 vccd1 _1756_/A sky130_fd_sc_hd__xnor2_2
XFILLER_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_i_clk clkbuf_4_9_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2806_/CLK sky130_fd_sc_hd__clkbuf_2
X_2205_ _2800_/Q _2657_/Q _2658_/Q _2204_/X vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__o31a_1
X_2136_ _2132_/X _2135_/Y _2132_/A _2070_/X vssd1 vssd1 vccd1 vccd1 _2739_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2067_ _2693_/Q vssd1 vssd1 vccd1 vccd1 _2068_/A sky130_fd_sc_hd__inv_2
XFILLER_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2754_ _2757_/CLK _2754_/D _2475_/Y vssd1 vssd1 vccd1 vccd1 _2754_/Q sky130_fd_sc_hd__dfrtp_1
X_1705_ _1713_/A _1713_/C vssd1 vssd1 vccd1 vccd1 _1737_/A sky130_fd_sc_hd__or2_1
X_2685_ _2726_/CLK _2685_/D vssd1 vssd1 vccd1 vccd1 _2685_/Q sky130_fd_sc_hd__dfxtp_1
X_1567_ _1581_/A _1576_/A _1581_/B _1595_/A _1566_/X vssd1 vssd1 vccd1 vccd1 _1577_/C
+ sky130_fd_sc_hd__a41o_1
X_1636_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1636_/Y sky130_fd_sc_hd__inv_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1498_ _1492_/X _1490_/Y _1496_/Y _1494_/A vssd1 vssd1 vccd1 vccd1 _1499_/B sky130_fd_sc_hd__a211o_1
X_2119_ _2113_/X _2117_/Y _2118_/X _2099_/X _2059_/A vssd1 vssd1 vccd1 vccd1 _2745_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1421_ _2752_/Q vssd1 vssd1 vccd1 vccd1 _2063_/A sky130_fd_sc_hd__clkbuf_2
X_2470_ _2470_/A vssd1 vssd1 vccd1 vccd1 _2475_/A sky130_fd_sc_hd__buf_2
X_1352_ _1352_/A vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__inv_2
X_2668_ _2760_/CLK _2668_/D vssd1 vssd1 vccd1 vccd1 _2668_/Q sky130_fd_sc_hd__dfxtp_1
X_2806_ _2806_/CLK _2806_/D vssd1 vssd1 vccd1 vccd1 _2806_/Q sky130_fd_sc_hd__dfxtp_1
X_2737_ _2759_/CLK _2737_/D _2455_/Y vssd1 vssd1 vccd1 vccd1 _2737_/Q sky130_fd_sc_hd__dfrtp_1
X_1619_ _1619_/A _1619_/B _1619_/C vssd1 vssd1 vccd1 vccd1 _1620_/B sky130_fd_sc_hd__and3_1
Xclkbuf_3_5_0_i_clk clkbuf_3_5_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_i_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_2599_ _2576_/X _2580_/Y _2590_/B _2598_/X _2797_/Q vssd1 vssd1 vccd1 vccd1 _2599_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1970_ _1978_/C vssd1 vssd1 vccd1 vccd1 _2026_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2522_ _2521_/X _2183_/B _2527_/A vssd1 vssd1 vccd1 vccd1 _2525_/B sky130_fd_sc_hd__o21ai_1
X_1404_ _1412_/A _1413_/S _1401_/X _1406_/A vssd1 vssd1 vccd1 vccd1 _1405_/B sky130_fd_sc_hd__o211a_1
X_2384_ _2386_/C _2384_/B vssd1 vssd1 vccd1 vccd1 _2702_/D sky130_fd_sc_hd__nor2_1
X_2453_ _2457_/A vssd1 vssd1 vccd1 vccd1 _2453_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1335_ _2735_/Q _2734_/Q _2733_/Q _2732_/Q vssd1 vssd1 vccd1 vccd1 _1510_/A sky130_fd_sc_hd__or4_1
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1953_ _1953_/A _1953_/B vssd1 vssd1 vccd1 vccd1 _1953_/Y sky130_fd_sc_hd__nand2_1
X_1884_ _1975_/A vssd1 vssd1 vccd1 vccd1 _1985_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2505_ _2781_/Q _2510_/C vssd1 vssd1 vccd1 vccd1 _2507_/C sky130_fd_sc_hd__or2_1
X_2298_ _2672_/Q _2298_/B vssd1 vssd1 vccd1 vccd1 _2300_/A sky130_fd_sc_hd__nor2_1
X_2436_ _2724_/Q _2435_/C _2725_/Q vssd1 vssd1 vccd1 vccd1 _2437_/B sky130_fd_sc_hd__a21oi_1
X_2367_ _2367_/A vssd1 vssd1 vccd1 vccd1 _2697_/D sky130_fd_sc_hd__clkbuf_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_i_clk clkbuf_2_3_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2221_ _2221_/A _2225_/B vssd1 vssd1 vccd1 vccd1 _2227_/C sky130_fd_sc_hd__or2_1
X_2152_ _2149_/B _2151_/Y _2053_/A _2070_/X vssd1 vssd1 vccd1 vccd1 _2734_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2083_ _2083_/A _2083_/B vssd1 vssd1 vccd1 vccd1 _2083_/X sky130_fd_sc_hd__or2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1936_ _1936_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1936_/X sky130_fd_sc_hd__or2_1
X_1867_ _1947_/A vssd1 vssd1 vccd1 vccd1 _1963_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_4_4_0_i_clk clkbuf_4_5_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2805_/CLK sky130_fd_sc_hd__clkbuf_2
X_1798_ _1798_/A _2006_/A vssd1 vssd1 vccd1 vccd1 _1910_/B sky130_fd_sc_hd__nor2_2
X_2419_ _2421_/C _2419_/B vssd1 vssd1 vccd1 vccd1 _2717_/D sky130_fd_sc_hd__nor2_1
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1721_ _1720_/Y _1720_/A _1721_/S vssd1 vssd1 vccd1 vccd1 _1743_/A sky130_fd_sc_hd__mux2_1
X_2770_ _2805_/CLK _2770_/D _2494_/Y vssd1 vssd1 vccd1 vccd1 _2770_/Q sky130_fd_sc_hd__dfrtp_2
X_1583_ _1595_/A _1620_/A _1585_/A _1619_/B _1587_/B vssd1 vssd1 vccd1 vccd1 _1591_/B
+ sky130_fd_sc_hd__a41o_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ _1901_/A _1661_/B vssd1 vssd1 vccd1 vccd1 _1665_/A sky130_fd_sc_hd__and2_2
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _2132_/A _2138_/A _2105_/X vssd1 vssd1 vccd1 vccd1 _2135_/Y sky130_fd_sc_hd__o21ai_1
X_2204_ _2804_/Q _2234_/B _2657_/D vssd1 vssd1 vccd1 vccd1 _2204_/X sky130_fd_sc_hd__a21o_1
X_2066_ _2757_/Q _2083_/A _2083_/B vssd1 vssd1 vccd1 vccd1 _2079_/A sky130_fd_sc_hd__and3_1
X_1919_ _1803_/X _1912_/A _1915_/B _1910_/B _1910_/A vssd1 vssd1 vccd1 vccd1 _1920_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2684_ _2726_/CLK _2684_/D vssd1 vssd1 vccd1 vccd1 _2684_/Q sky130_fd_sc_hd__dfxtp_1
X_2753_ _2757_/CLK _2753_/D _2474_/Y vssd1 vssd1 vccd1 vccd1 _2753_/Q sky130_fd_sc_hd__dfrtp_1
X_1704_ _1704_/A _1704_/B vssd1 vssd1 vccd1 vccd1 _1713_/A sky130_fd_sc_hd__or2_1
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1566_ _1555_/A _1565_/Y _1578_/B vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__o21a_1
X_1635_ _1900_/A _1635_/B vssd1 vssd1 vccd1 vccd1 _1636_/A sky130_fd_sc_hd__or2_1
X_1497_ _1494_/A _1492_/X _1496_/Y vssd1 vssd1 vccd1 vccd1 _1499_/A sky130_fd_sc_hd__o21ai_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2118_ _2121_/A _2058_/A _2126_/A _2059_/A vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__a31o_1
X_2049_ _2741_/Q vssd1 vssd1 vccd1 vccd1 _2130_/A sky130_fd_sc_hd__clkbuf_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_i_clk clkbuf_3_1_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1420_ _1420_/A vssd1 vssd1 vccd1 vccd1 _1551_/B sky130_fd_sc_hd__clkbuf_2
X_1351_ _2747_/Q _1351_/B vssd1 vssd1 vccd1 vccd1 _1352_/A sky130_fd_sc_hd__xnor2_2
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2805_ _2805_/CLK _2805_/D vssd1 vssd1 vccd1 vccd1 _2805_/Q sky130_fd_sc_hd__dfxtp_2
X_1618_ _1618_/A _1618_/B vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__or2_1
X_2667_ _2673_/CLK _2667_/D vssd1 vssd1 vccd1 vccd1 _2667_/Q sky130_fd_sc_hd__dfxtp_1
X_2736_ _2759_/CLK _2736_/D _2454_/Y vssd1 vssd1 vccd1 vccd1 _2736_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1549_ _1549_/A _1549_/B vssd1 vssd1 vccd1 vccd1 _1563_/A sky130_fd_sc_hd__and2_1
X_2598_ _2598_/A vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2521_ _2622_/C vssd1 vssd1 vccd1 vccd1 _2521_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1403_ _1403_/A _1407_/B vssd1 vssd1 vccd1 vccd1 _1413_/S sky130_fd_sc_hd__xnor2_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1334_ _1334_/A vssd1 vssd1 vccd1 vccd1 _1512_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2383_ _2702_/Q _2383_/B vssd1 vssd1 vccd1 vccd1 _2384_/B sky130_fd_sc_hd__nor2_1
X_2452_ _2470_/A vssd1 vssd1 vccd1 vccd1 _2457_/A sky130_fd_sc_hd__buf_2
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2719_ _2807_/CLK _2719_/D vssd1 vssd1 vccd1 vccd1 _2719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1952_ _1935_/B _2013_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1953_/B sky130_fd_sc_hd__o21ai_1
X_1883_ _1883_/A _1883_/B vssd1 vssd1 vccd1 vccd1 _1975_/A sky130_fd_sc_hd__nor2_1
X_2435_ _2725_/Q _2724_/Q _2435_/C vssd1 vssd1 vccd1 vccd1 _2439_/B sky130_fd_sc_hd__and3_1
X_2504_ _2780_/Q _2502_/B _2503_/Y vssd1 vssd1 vccd1 vccd1 _2780_/D sky130_fd_sc_hd__o21a_1
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2297_ _2297_/A _2298_/B vssd1 vssd1 vccd1 vccd1 _2671_/D sky130_fd_sc_hd__nor2_1
X_2366_ _2380_/A _2366_/B _2366_/C vssd1 vssd1 vccd1 vccd1 _2367_/A sky130_fd_sc_hd__and3_1
Xclkbuf_4_0_0_i_clk clkbuf_4_1_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2783_/CLK sky130_fd_sc_hd__clkbuf_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2220_ _2221_/A _2225_/B vssd1 vssd1 vccd1 vccd1 _2222_/B sky130_fd_sc_hd__nand2_1
X_2082_ _2083_/A _2083_/B vssd1 vssd1 vccd1 vccd1 _2082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2151_ _2053_/A _2154_/A _2113_/A vssd1 vssd1 vccd1 vccd1 _2151_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1935_ _1936_/B _1935_/B _1935_/C vssd1 vssd1 vccd1 vccd1 _1953_/A sky130_fd_sc_hd__or3_1
X_1866_ _1877_/A _1878_/A vssd1 vssd1 vccd1 vccd1 _1866_/X sky130_fd_sc_hd__and2_1
X_1797_ _1817_/B vssd1 vssd1 vccd1 vccd1 _1798_/A sky130_fd_sc_hd__inv_2
X_2418_ _2717_/Q _2418_/B vssd1 vssd1 vccd1 vccd1 _2419_/B sky130_fd_sc_hd__nor2_1
X_2349_ _2349_/A _2349_/B _2349_/C vssd1 vssd1 vccd1 vccd1 _2356_/B sky130_fd_sc_hd__or3_1
XFILLER_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1651_ _1900_/A _1651_/B vssd1 vssd1 vccd1 vccd1 _1661_/B sky130_fd_sc_hd__xor2_1
X_1720_ _1720_/A _1720_/B vssd1 vssd1 vccd1 vccd1 _1720_/Y sky130_fd_sc_hd__nand2_1
X_1582_ _1577_/X _1580_/X _1581_/Y vssd1 vssd1 vccd1 vccd1 _1587_/B sky130_fd_sc_hd__o21a_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2065_ _2065_/A _2089_/A vssd1 vssd1 vccd1 vccd1 _2083_/B sky130_fd_sc_hd__and2_1
X_2134_ _2130_/B _2133_/Y _2056_/A _2070_/X vssd1 vssd1 vccd1 vccd1 _2740_/D sky130_fd_sc_hd__a2bb2o_1
X_2203_ _2805_/Q _2657_/D _2200_/X _2202_/X vssd1 vssd1 vccd1 vccd1 _2227_/A sky130_fd_sc_hd__o211a_1
X_1918_ _1918_/A _1918_/B vssd1 vssd1 vccd1 vccd1 _1930_/B sky130_fd_sc_hd__xor2_1
X_1849_ _1857_/A _1849_/B vssd1 vssd1 vccd1 vccd1 _1862_/A sky130_fd_sc_hd__and2_1
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2683_ _2726_/CLK _2683_/D vssd1 vssd1 vccd1 vccd1 _2683_/Q sky130_fd_sc_hd__dfxtp_1
X_1634_ _1642_/A _1642_/B vssd1 vssd1 vccd1 vccd1 _1635_/B sky130_fd_sc_hd__xnor2_1
X_2752_ _2757_/CLK _2752_/D _2473_/Y vssd1 vssd1 vccd1 vccd1 _2752_/Q sky130_fd_sc_hd__dfrtp_1
X_1703_ _1739_/A vssd1 vssd1 vccd1 vccd1 _1703_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1565_ _1578_/A _1897_/C _1565_/C vssd1 vssd1 vccd1 vccd1 _1565_/Y sky130_fd_sc_hd__nor3_1
X_1496_ _1496_/A _1496_/B vssd1 vssd1 vccd1 vccd1 _1496_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2117_ _2117_/A vssd1 vssd1 vccd1 vccd1 _2117_/Y sky130_fd_sc_hd__inv_2
X_2048_ _2744_/Q vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1350_ _1512_/A _2746_/Q _1348_/B vssd1 vssd1 vccd1 vccd1 _1351_/B sky130_fd_sc_hd__a21bo_1
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2804_ _2809_/CLK _2804_/D vssd1 vssd1 vccd1 vccd1 _2804_/Q sky130_fd_sc_hd__dfxtp_2
X_1617_ _1603_/Y _1604_/Y _1630_/A _1611_/Y _1637_/A vssd1 vssd1 vccd1 vccd1 _1624_/B
+ sky130_fd_sc_hd__a2111o_1
X_2666_ _2673_/CLK _2666_/D vssd1 vssd1 vccd1 vccd1 _2666_/Q sky130_fd_sc_hd__dfxtp_1
X_2597_ _2576_/X _2577_/X _2618_/A vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__a21o_1
X_2735_ _2759_/CLK _2735_/D _2453_/Y vssd1 vssd1 vccd1 vccd1 _2735_/Q sky130_fd_sc_hd__dfrtp_1
X_1548_ _1590_/A _1590_/B vssd1 vssd1 vccd1 vccd1 _1899_/A sky130_fd_sc_hd__or2_2
X_1479_ _1479_/A _1479_/B vssd1 vssd1 vccd1 vccd1 _1483_/B sky130_fd_sc_hd__or2_1
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1402_ _1406_/A _1412_/A _1401_/X vssd1 vssd1 vccd1 vccd1 _1405_/A sky130_fd_sc_hd__a21oi_1
X_2520_ _2786_/Q vssd1 vssd1 vccd1 vccd1 _2622_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_2451_ _2451_/A vssd1 vssd1 vccd1 vccd1 _2451_/Y sky130_fd_sc_hd__inv_2
X_1333_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2382_ _2701_/Q _2702_/Q _2382_/C vssd1 vssd1 vccd1 vccd1 _2386_/C sky130_fd_sc_hd__and3_1
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2718_ _2807_/CLK _2718_/D vssd1 vssd1 vccd1 vccd1 _2718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2649_ _2807_/Q _2655_/B _2648_/X _2636_/X vssd1 vssd1 vccd1 vccd1 _2807_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1951_ _1951_/A _1951_/B vssd1 vssd1 vccd1 vccd1 _1951_/Y sky130_fd_sc_hd__nand2_1
X_1882_ _1883_/A _1883_/B _1875_/A vssd1 vssd1 vccd1 vccd1 _1890_/B sky130_fd_sc_hd__o21a_1
X_2434_ _2724_/Q _2435_/C vssd1 vssd1 vccd1 vccd1 _2724_/D sky130_fd_sc_hd__xor2_1
X_2365_ _2697_/Q _2696_/Q vssd1 vssd1 vccd1 vccd1 _2366_/C sky130_fd_sc_hd__nand2_1
X_2503_ _2503_/A _2510_/C vssd1 vssd1 vccd1 vccd1 _2503_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2296_ _2671_/Q _2299_/C vssd1 vssd1 vccd1 vccd1 _2298_/B sky130_fd_sc_hd__and2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2081_ _2073_/X _2079_/Y _2080_/X _2077_/X _2757_/Q vssd1 vssd1 vccd1 vccd1 _2757_/D
+ sky130_fd_sc_hd__a32o_1
X_2150_ _2137_/X _2148_/Y _2149_/X _2146_/X _2149_/A vssd1 vssd1 vccd1 vccd1 _2735_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1934_ _1803_/X _1913_/B _1933_/X vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__a21bo_1
X_1865_ _1870_/B _1947_/A vssd1 vssd1 vccd1 vccd1 _1878_/A sky130_fd_sc_hd__xor2_1
X_1796_ _1801_/B vssd1 vssd1 vccd1 vccd1 _2006_/A sky130_fd_sc_hd__buf_2
X_2348_ _2725_/Q _2724_/Q _2727_/Q _2726_/Q vssd1 vssd1 vccd1 vccd1 _2349_/C sky130_fd_sc_hd__or4_1
X_2417_ _2717_/Q _2418_/B vssd1 vssd1 vccd1 vccd1 _2421_/C sky130_fd_sc_hd__and2_1
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2279_ _2285_/A _2279_/B _2279_/C vssd1 vssd1 vccd1 vccd1 _2280_/A sky130_fd_sc_hd__and3_1
XFILLER_52_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1581_ _1581_/A _1581_/B _1581_/C vssd1 vssd1 vccd1 vccd1 _1581_/Y sky130_fd_sc_hd__nand3_1
X_1650_ _1636_/Y _1640_/X _1649_/X vssd1 vssd1 vccd1 vccd1 _1650_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_7_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2809_/Q _2657_/D _2234_/B vssd1 vssd1 vccd1 vccd1 _2202_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2064_ _2064_/A _2093_/A _2093_/B vssd1 vssd1 vccd1 vccd1 _2089_/A sky130_fd_sc_hd__and3_1
X_2133_ _2056_/A _2132_/X _2105_/X vssd1 vssd1 vccd1 vccd1 _2133_/Y sky130_fd_sc_hd__o21ai_1
X_1917_ _1917_/A _1914_/A vssd1 vssd1 vccd1 vccd1 _1918_/B sky130_fd_sc_hd__or2b_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1848_ _1851_/A _1850_/A vssd1 vssd1 vccd1 vccd1 _1849_/B sky130_fd_sc_hd__xor2_1
X_1779_ _1811_/A vssd1 vssd1 vccd1 vccd1 _1779_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2751_ _2758_/CLK _2751_/D _2472_/Y vssd1 vssd1 vccd1 vccd1 _2751_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1564_ _1564_/A _1570_/A _1570_/B _1571_/A vssd1 vssd1 vccd1 vccd1 _1581_/B sky130_fd_sc_hd__or4b_2
X_1633_ _1638_/A _1638_/B _1629_/X _1632_/X vssd1 vssd1 vccd1 vccd1 _1642_/B sky130_fd_sc_hd__o31ai_4
X_2682_ _2726_/CLK _2682_/D vssd1 vssd1 vccd1 vccd1 _2682_/Q sky130_fd_sc_hd__dfxtp_1
X_1702_ _1720_/A _1721_/S _1720_/B vssd1 vssd1 vccd1 vccd1 _1731_/A sky130_fd_sc_hd__a21oi_4
X_1495_ _1546_/A _1546_/B _1483_/A vssd1 vssd1 vccd1 vccd1 _1496_/A sky130_fd_sc_hd__a21oi_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ _2746_/Q vssd1 vssd1 vccd1 vccd1 _2115_/A sky130_fd_sc_hd__clkbuf_1
X_2116_ _2113_/X _2114_/Y _2115_/X _2099_/X _2115_/A vssd1 vssd1 vccd1 vccd1 _2746_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2803_ _2805_/CLK _2803_/D vssd1 vssd1 vccd1 vccd1 _2803_/Q sky130_fd_sc_hd__dfxtp_1
X_2734_ _2759_/CLK _2734_/D _2451_/Y vssd1 vssd1 vccd1 vccd1 _2734_/Q sky130_fd_sc_hd__dfrtp_1
X_2665_ _2760_/CLK _2665_/D vssd1 vssd1 vccd1 vccd1 _2665_/Q sky130_fd_sc_hd__dfxtp_1
X_1616_ _1618_/B _1616_/B vssd1 vssd1 vccd1 vccd1 _1637_/A sky130_fd_sc_hd__nand2_1
X_1547_ _1899_/C vssd1 vssd1 vccd1 vccd1 _1642_/A sky130_fd_sc_hd__inv_2
X_2596_ _2600_/A _2600_/B vssd1 vssd1 vccd1 vccd1 _2618_/A sky130_fd_sc_hd__nand2_1
X_1478_ _1485_/B _1485_/C _1471_/X _1485_/A vssd1 vssd1 vccd1 vccd1 _1479_/B sky130_fd_sc_hd__a211oi_1
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1401_ _1407_/B _1407_/C vssd1 vssd1 vccd1 vccd1 _1401_/X sky130_fd_sc_hd__or2_1
X_2381_ _2381_/A vssd1 vssd1 vccd1 vccd1 _2701_/D sky130_fd_sc_hd__clkbuf_1
X_2450_ _2451_/A vssd1 vssd1 vccd1 vccd1 _2450_/Y sky130_fd_sc_hd__inv_2
X_1332_ _1373_/A vssd1 vssd1 vccd1 vccd1 _1410_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2717_ _2727_/CLK _2717_/D vssd1 vssd1 vccd1 vccd1 _2717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2648_ _2807_/Q _2242_/A _2183_/Y _2625_/A _2647_/X vssd1 vssd1 vccd1 vccd1 _2648_/X
+ sky130_fd_sc_hd__a311o_1
X_2579_ _2805_/Q _2632_/B _2578_/X _2183_/A vssd1 vssd1 vccd1 vccd1 _2593_/A sky130_fd_sc_hd__a22o_1
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1950_ _1948_/Y _1937_/X _1949_/X vssd1 vssd1 vccd1 vccd1 _1965_/C sky130_fd_sc_hd__a21o_1
X_2502_ _2780_/Q _2502_/B vssd1 vssd1 vccd1 vccd1 _2510_/C sky130_fd_sc_hd__and2_1
X_1881_ _1869_/Y _1976_/A _1880_/X vssd1 vssd1 vccd1 vccd1 _1883_/B sky130_fd_sc_hd__o21ai_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2433_ _2435_/C _2433_/B vssd1 vssd1 vccd1 vccd1 _2723_/D sky130_fd_sc_hd__nor2_1
X_2364_ _2697_/Q _2696_/Q vssd1 vssd1 vccd1 vccd1 _2366_/B sky130_fd_sc_hd__or2_1
X_2295_ _2671_/Q _2299_/C vssd1 vssd1 vccd1 vccd1 _2297_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2810__27 vssd1 vssd1 vccd1 vccd1 o_display_cathode[7] _2810__27/LO sky130_fd_sc_hd__conb_1
XFILLER_11_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ _2083_/A _2065_/A _2089_/A _2757_/Q vssd1 vssd1 vccd1 vccd1 _2080_/X sky130_fd_sc_hd__a31o_1
XFILLER_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1933_ _1913_/A _1912_/A _1915_/B _1803_/A vssd1 vssd1 vccd1 vccd1 _1933_/X sky130_fd_sc_hd__a31o_1
X_1864_ _1858_/X _1872_/S _1863_/X vssd1 vssd1 vccd1 vccd1 _1947_/A sky130_fd_sc_hd__o21ai_2
X_1795_ _1819_/S _1910_/A _1817_/B _1920_/A _1818_/B vssd1 vssd1 vccd1 vccd1 _1801_/B
+ sky130_fd_sc_hd__a41oi_1
X_2278_ _2284_/C vssd1 vssd1 vccd1 vccd1 _2279_/C sky130_fd_sc_hd__clkinv_2
X_2347_ _2713_/Q _2712_/Q _2715_/Q _2714_/Q vssd1 vssd1 vccd1 vccd1 _2349_/B sky130_fd_sc_hd__or4_1
X_2416_ _2418_/B _2416_/B vssd1 vssd1 vccd1 vccd1 _2716_/D sky130_fd_sc_hd__nor2_1
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1580_ _1897_/C _1565_/C _1578_/X _1579_/X _1581_/A vssd1 vssd1 vccd1 vccd1 _1580_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2658_/Q vssd1 vssd1 vccd1 vccd1 _2234_/B sky130_fd_sc_hd__clkinv_2
X_2132_ _2132_/A _2138_/A vssd1 vssd1 vccd1 vccd1 _2132_/X sky130_fd_sc_hd__and2_1
X_2063_ _2063_/A _2097_/A vssd1 vssd1 vccd1 vccd1 _2093_/B sky130_fd_sc_hd__and2_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1916_ _1928_/A _1929_/A vssd1 vssd1 vccd1 vccd1 _1930_/A sky130_fd_sc_hd__nor2_1
X_1847_ _1847_/A _1847_/B vssd1 vssd1 vccd1 vccd1 _1850_/A sky130_fd_sc_hd__or2_1
X_1778_ _1778_/A _1807_/A vssd1 vssd1 vccd1 vccd1 _1811_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2681_ _2726_/CLK _2681_/D vssd1 vssd1 vccd1 vccd1 _2681_/Q sky130_fd_sc_hd__dfxtp_1
X_2750_ _2758_/CLK _2750_/D _2471_/Y vssd1 vssd1 vccd1 vccd1 _2750_/Q sky130_fd_sc_hd__dfrtp_2
X_1701_ _1537_/X _1538_/Y _1700_/X vssd1 vssd1 vccd1 vccd1 _1720_/B sky130_fd_sc_hd__a21boi_2
XFILLER_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1632_ _1611_/Y _1631_/X _1624_/B vssd1 vssd1 vccd1 vccd1 _1632_/X sky130_fd_sc_hd__a21bo_1
X_1563_ _1563_/A _1563_/B _1578_/B vssd1 vssd1 vccd1 vccd1 _1570_/B sky130_fd_sc_hd__and3_1
X_1494_ _1494_/A _1501_/A vssd1 vssd1 vccd1 vccd1 _1519_/A sky130_fd_sc_hd__xnor2_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2115_ _2115_/A _2117_/A vssd1 vssd1 vccd1 vccd1 _2115_/X sky130_fd_sc_hd__or2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ _2750_/Q vssd1 vssd1 vccd1 vccd1 _2102_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2664_ _2760_/CLK _2664_/D vssd1 vssd1 vccd1 vccd1 _2664_/Q sky130_fd_sc_hd__dfxtp_1
X_2733_ _2759_/CLK _2733_/D _2450_/Y vssd1 vssd1 vccd1 vccd1 _2733_/Q sky130_fd_sc_hd__dfrtp_1
X_2802_ _2802_/CLK _2802_/D vssd1 vssd1 vccd1 vccd1 _2802_/Q sky130_fd_sc_hd__dfxtp_1
X_1615_ _1612_/Y _1613_/X _1614_/Y vssd1 vssd1 vccd1 vccd1 _1616_/B sky130_fd_sc_hd__a21o_1
X_1477_ _1477_/A _1477_/B vssd1 vssd1 vccd1 vccd1 _1485_/C sky130_fd_sc_hd__or2_1
X_1546_ _1546_/A _1546_/B vssd1 vssd1 vccd1 vccd1 _1899_/C sky130_fd_sc_hd__nand2_1
X_2595_ _2777_/Q _2190_/X _2554_/A vssd1 vssd1 vccd1 vccd1 _2600_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2029_ _2029_/A _2029_/B vssd1 vssd1 vccd1 vccd1 _2034_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1400_ _1393_/Y _1553_/A _1553_/B vssd1 vssd1 vccd1 vccd1 _1407_/C sky130_fd_sc_hd__and3b_1
X_1331_ _2759_/Q vssd1 vssd1 vccd1 vccd1 _1373_/A sky130_fd_sc_hd__clkbuf_2
X_2380_ _2380_/A _2380_/B _2380_/C vssd1 vssd1 vccd1 vccd1 _2381_/A sky130_fd_sc_hd__and3_1
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2716_ _2807_/CLK _2716_/D vssd1 vssd1 vccd1 vccd1 _2716_/Q sky130_fd_sc_hd__dfxtp_1
X_2647_ _2242_/A _2195_/X _2605_/Y _2248_/A _2806_/Q vssd1 vssd1 vccd1 vccd1 _2647_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1529_ _1529_/A _1529_/B vssd1 vssd1 vccd1 vccd1 _1529_/X sky130_fd_sc_hd__or2_1
X_2578_ _2801_/Q _2809_/Q _2581_/A vssd1 vssd1 vccd1 vccd1 _2578_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2822__25 vssd1 vssd1 vccd1 vccd1 _2822__25/HI o_io_oeb[11] sky130_fd_sc_hd__conb_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1870_/A _1866_/X _1872_/X vssd1 vssd1 vccd1 vccd1 _1880_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2501_ _2779_/Q _2497_/B _2500_/Y vssd1 vssd1 vccd1 vccd1 _2779_/D sky130_fd_sc_hd__o21a_1
X_2294_ _2294_/A _2299_/C vssd1 vssd1 vccd1 vccd1 _2670_/D sky130_fd_sc_hd__nor2_1
X_2432_ _2723_/Q _2432_/B vssd1 vssd1 vccd1 vccd1 _2433_/B sky130_fd_sc_hd__nor2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2363_ _2444_/A vssd1 vssd1 vccd1 vccd1 _2363_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1932_ _1935_/B _2013_/A _1931_/Y vssd1 vssd1 vccd1 vccd1 _1951_/B sky130_fd_sc_hd__o21a_1
X_1863_ _1853_/B _1862_/X _1856_/A vssd1 vssd1 vccd1 vccd1 _1863_/X sky130_fd_sc_hd__a21o_1
X_2415_ _2715_/Q _2414_/C _2716_/Q vssd1 vssd1 vccd1 vccd1 _2416_/B sky130_fd_sc_hd__a21oi_1
X_1794_ _1791_/X _1792_/Y _1794_/S vssd1 vssd1 vccd1 vccd1 _1818_/B sky130_fd_sc_hd__mux2_1
X_2277_ _2664_/Q _2663_/Q _2665_/Q _2277_/D vssd1 vssd1 vccd1 vccd1 _2284_/C sky130_fd_sc_hd__and4_1
X_2346_ _2717_/Q _2716_/Q _2719_/Q _2718_/Q vssd1 vssd1 vccd1 vccd1 _2349_/A sky130_fd_sc_hd__or4_1
XFILLER_37_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2062_ _2751_/Q _2102_/A _2102_/B vssd1 vssd1 vccd1 vccd1 _2097_/A sky130_fd_sc_hd__and3_1
X_2131_ _2113_/X _2129_/Y _2130_/X _2122_/X _2130_/A vssd1 vssd1 vccd1 vccd1 _2741_/D
+ sky130_fd_sc_hd__a32o_1
X_2200_ _2801_/Q _2657_/Q _2658_/Q vssd1 vssd1 vccd1 vccd1 _2200_/X sky130_fd_sc_hd__or3_1
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1915_ _1917_/A _1915_/B vssd1 vssd1 vccd1 vccd1 _1929_/A sky130_fd_sc_hd__xor2_2
X_1846_ _1810_/X _1917_/A _1845_/X vssd1 vssd1 vccd1 vccd1 _1847_/B sky130_fd_sc_hd__o21ai_1
X_1777_ _2055_/B _1777_/B vssd1 vssd1 vccd1 vccd1 _1807_/A sky130_fd_sc_hd__xnor2_2
XFILLER_57_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2329_ _2329_/A _2332_/C vssd1 vssd1 vccd1 vccd1 _2684_/D sky130_fd_sc_hd__nor2_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1631_ _1611_/Y _1624_/C _1630_/X _1626_/Y vssd1 vssd1 vccd1 vccd1 _1631_/X sky130_fd_sc_hd__a211o_1
X_2680_ _2726_/CLK _2680_/D vssd1 vssd1 vccd1 vccd1 _2680_/Q sky130_fd_sc_hd__dfxtp_1
X_1700_ _1537_/X _1541_/X _1538_/Y vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__a21o_1
X_1562_ _1431_/C _1563_/B _1441_/X vssd1 vssd1 vccd1 vccd1 _1564_/A sky130_fd_sc_hd__o21ai_1
X_1493_ _1488_/X _1490_/Y _1492_/X vssd1 vssd1 vccd1 vccd1 _1501_/A sky130_fd_sc_hd__o21ai_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2114_ _2115_/A _2117_/A vssd1 vssd1 vccd1 vccd1 _2114_/Y sky130_fd_sc_hd__nand2_1
X_2045_ _2753_/Q vssd1 vssd1 vccd1 vccd1 _2093_/A sky130_fd_sc_hd__clkbuf_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1829_ _2157_/A _1829_/B vssd1 vssd1 vccd1 vccd1 _1829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2801_ _2809_/CLK _2801_/D vssd1 vssd1 vccd1 vccd1 _2801_/Q sky130_fd_sc_hd__dfxtp_1
X_2663_ _2760_/CLK _2663_/D vssd1 vssd1 vccd1 vccd1 _2663_/Q sky130_fd_sc_hd__dfxtp_1
X_1614_ _1614_/A _1614_/B vssd1 vssd1 vccd1 vccd1 _1614_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2732_ _2759_/CLK _2732_/D _2449_/Y vssd1 vssd1 vccd1 vccd1 _2732_/Q sky130_fd_sc_hd__dfrtp_1
X_2594_ _2577_/A _2621_/A _2777_/Q vssd1 vssd1 vccd1 vccd1 _2600_/A sky130_fd_sc_hd__o21ai_1
X_1476_ _1470_/A _1590_/B _1474_/Y vssd1 vssd1 vccd1 vccd1 _1477_/B sky130_fd_sc_hd__a21oi_1
X_1545_ _1545_/A _1545_/B vssd1 vssd1 vccd1 vccd1 _1901_/A sky130_fd_sc_hd__and2_1
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2028_ _2028_/A vssd1 vssd1 vccd1 vccd1 _2763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1330_ _1326_/Y _2692_/D _2694_/D _2770_/Q vssd1 vssd1 vccd1 vccd1 _2770_/D sky130_fd_sc_hd__o22a_1
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2715_ _2727_/CLK _2715_/D vssd1 vssd1 vccd1 vccd1 _2715_/Q sky130_fd_sc_hd__dfxtp_1
X_2646_ _2646_/A vssd1 vssd1 vccd1 vccd1 _2806_/D sky130_fd_sc_hd__clkbuf_1
X_2577_ _2577_/A _2622_/A _2622_/C vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__or3_1
X_1459_ _1462_/A _1461_/A _1457_/Y _1458_/X vssd1 vssd1 vccd1 vccd1 _1470_/B sky130_fd_sc_hd__o2bb2a_1
X_1528_ _1530_/A _1901_/B _1527_/A vssd1 vssd1 vccd1 vccd1 _1529_/B sky130_fd_sc_hd__o21a_1
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2431_ _2723_/Q _2432_/B vssd1 vssd1 vccd1 vccd1 _2435_/C sky130_fd_sc_hd__and2_1
X_2500_ _2503_/A _2502_/B vssd1 vssd1 vccd1 vccd1 _2500_/Y sky130_fd_sc_hd__nor2_1
X_2293_ _2670_/Q _2669_/Q _2293_/C vssd1 vssd1 vccd1 vccd1 _2299_/C sky130_fd_sc_hd__and3_1
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2362_ _2444_/A vssd1 vssd1 vccd1 vccd1 _2362_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2629_ _2803_/Q _2605_/Y _2629_/S vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1931_ _1930_/A _1920_/Y _1930_/B vssd1 vssd1 vccd1 vccd1 _1931_/Y sky130_fd_sc_hd__o21ai_1
X_1862_ _1862_/A _1856_/B vssd1 vssd1 vccd1 vccd1 _1862_/X sky130_fd_sc_hd__or2b_1
X_1793_ _1793_/A _1793_/B _1793_/C _1793_/D vssd1 vssd1 vccd1 vccd1 _1794_/S sky130_fd_sc_hd__and4_1
X_2414_ _2715_/Q _2716_/Q _2414_/C vssd1 vssd1 vccd1 vccd1 _2418_/B sky130_fd_sc_hd__and3_1
X_2276_ _2664_/Q _2663_/Q _2262_/A _2665_/Q vssd1 vssd1 vccd1 vccd1 _2279_/B sky130_fd_sc_hd__a31o_1
X_2345_ _2721_/Q _2720_/Q _2723_/Q _2722_/Q vssd1 vssd1 vccd1 vccd1 _2356_/A sky130_fd_sc_hd__or4_1
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2061_ _2749_/Q _2104_/A _2110_/A vssd1 vssd1 vccd1 vccd1 _2102_/B sky130_fd_sc_hd__and3_1
X_2130_ _2130_/A _2130_/B vssd1 vssd1 vccd1 vccd1 _2130_/X sky130_fd_sc_hd__or2_1
XFILLER_19_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1914_ _1914_/A vssd1 vssd1 vccd1 vccd1 _1915_/B sky130_fd_sc_hd__buf_2
X_1845_ _1778_/A _1808_/X _1812_/X vssd1 vssd1 vccd1 vccd1 _1845_/X sky130_fd_sc_hd__a21o_1
X_1776_ _1776_/A _1786_/A vssd1 vssd1 vccd1 vccd1 _1778_/A sky130_fd_sc_hd__xnor2_1
X_2328_ _2684_/Q _2328_/B vssd1 vssd1 vccd1 vccd1 _2332_/C sky130_fd_sc_hd__and2_1
X_2259_ _2262_/A _2259_/B vssd1 vssd1 vccd1 vccd1 _2662_/D sky130_fd_sc_hd__nor2_1
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1630_ _1630_/A _1637_/A vssd1 vssd1 vccd1 vccd1 _1630_/X sky130_fd_sc_hd__or2_1
X_1561_ _1561_/A _1570_/A vssd1 vssd1 vccd1 vccd1 _1576_/A sky130_fd_sc_hd__xnor2_2
X_1492_ _1483_/B _1491_/X _1546_/A vssd1 vssd1 vccd1 vccd1 _1492_/X sky130_fd_sc_hd__a21bo_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ _2113_/A vssd1 vssd1 vccd1 vccd1 _2113_/X sky130_fd_sc_hd__clkbuf_2
X_2044_ _2756_/Q vssd1 vssd1 vccd1 vccd1 _2083_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1828_ _2052_/B vssd1 vssd1 vccd1 vccd1 _2157_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1759_ _1754_/X _1755_/Y _1758_/X vssd1 vssd1 vccd1 vccd1 _1903_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2800_ _2806_/CLK _2800_/D vssd1 vssd1 vccd1 vccd1 _2800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2731_ _2802_/CLK _2731_/D _2448_/Y vssd1 vssd1 vccd1 vccd1 _2731_/Q sky130_fd_sc_hd__dfrtp_4
X_2662_ _2673_/CLK _2662_/D vssd1 vssd1 vccd1 vccd1 _2662_/Q sky130_fd_sc_hd__dfxtp_1
X_1613_ _1599_/A _1613_/B vssd1 vssd1 vccd1 vccd1 _1613_/X sky130_fd_sc_hd__and2b_1
X_1544_ _1544_/A vssd1 vssd1 vccd1 vccd1 _1672_/A sky130_fd_sc_hd__inv_2
X_2593_ _2593_/A _2611_/A vssd1 vssd1 vccd1 vccd1 _2621_/A sky130_fd_sc_hd__nor2_1
X_1475_ _1590_/A _1470_/C _1474_/Y _1470_/A vssd1 vssd1 vccd1 vccd1 _1477_/A sky130_fd_sc_hd__o211a_1
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2027_ _2763_/Q _2026_/Y _2032_/S vssd1 vssd1 vccd1 vccd1 _2028_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2714_ _2760_/CLK _2714_/D vssd1 vssd1 vccd1 vccd1 _2714_/Q sky130_fd_sc_hd__dfxtp_1
X_1527_ _1527_/A _1530_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1529_/A sky130_fd_sc_hd__nor3_1
X_2645_ _2645_/A _2645_/B vssd1 vssd1 vccd1 vccd1 _2646_/A sky130_fd_sc_hd__and2_1
X_2576_ _2576_/A vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1458_ _1458_/A _1458_/B _1591_/A vssd1 vssd1 vccd1 vccd1 _1458_/X sky130_fd_sc_hd__and3_1
X_1389_ _1383_/B _1383_/C _1555_/A _1388_/Y vssd1 vssd1 vccd1 vccd1 _1391_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2813__16 vssd1 vssd1 vccd1 vccd1 _2813__16/HI o_io_oeb[2] sky130_fd_sc_hd__conb_1
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2430_ _2432_/B _2430_/B vssd1 vssd1 vccd1 vccd1 _2722_/D sky130_fd_sc_hd__nor2_1
X_2361_ _2444_/A vssd1 vssd1 vccd1 vccd1 _2361_/Y sky130_fd_sc_hd__inv_2
X_2292_ _2669_/Q _2293_/C _2670_/Q vssd1 vssd1 vccd1 vccd1 _2294_/A sky130_fd_sc_hd__a21oi_1
XFILLER_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2559_ _2766_/Q _2793_/Q _2598_/A vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__mux2_1
X_2628_ _2802_/Q _2617_/X _2627_/X _2358_/X vssd1 vssd1 vccd1 vccd1 _2802_/D sky130_fd_sc_hd__o211a_1
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1930_ _1930_/A _1930_/B vssd1 vssd1 vccd1 vccd1 _1935_/B sky130_fd_sc_hd__or2_1
X_1861_ _1862_/A _1856_/B _1860_/Y vssd1 vssd1 vccd1 vccd1 _1872_/S sky130_fd_sc_hd__a21oi_1
X_1792_ _1792_/A vssd1 vssd1 vccd1 vccd1 _1792_/Y sky130_fd_sc_hd__clkinv_2
X_2344_ _2690_/Q _2342_/Y _2343_/Y _2689_/Q vssd1 vssd1 vccd1 vccd1 _2690_/D sky130_fd_sc_hd__a22o_1
X_2413_ _2715_/Q _2414_/C vssd1 vssd1 vccd1 vccd1 _2715_/D sky130_fd_sc_hd__xor2_1
X_2275_ _2664_/Q _2275_/B vssd1 vssd1 vccd1 vccd1 _2664_/D sky130_fd_sc_hd__xnor2_1
XFILLER_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _2747_/Q _2115_/A _2117_/A vssd1 vssd1 vccd1 vccd1 _2110_/A sky130_fd_sc_hd__and3_1
X_1913_ _1913_/A _1913_/B vssd1 vssd1 vccd1 vccd1 _1924_/A sky130_fd_sc_hd__xnor2_1
XFILLER_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1844_ _1854_/B _1854_/A vssd1 vssd1 vccd1 vccd1 _1847_/A sky130_fd_sc_hd__and2b_1
X_1775_ _1775_/A _1775_/B vssd1 vssd1 vccd1 vccd1 _1910_/A sky130_fd_sc_hd__xnor2_4
X_2258_ _2662_/Q _2258_/B vssd1 vssd1 vccd1 vccd1 _2259_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2327_ _2684_/Q _2328_/B vssd1 vssd1 vccd1 vccd1 _2329_/A sky130_fd_sc_hd__nor2_1
X_2189_ _2445_/A vssd1 vssd1 vccd1 vccd1 _2489_/A sky130_fd_sc_hd__buf_2
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1560_ _1578_/A _1578_/B _1563_/B vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__a21oi_2
Xclkbuf_4_13_0_i_clk clkbuf_3_6_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _2758_/CLK sky130_fd_sc_hd__clkbuf_2
X_1491_ _1490_/A _1349_/A _1483_/B _1546_/B vssd1 vssd1 vccd1 vccd1 _1491_/X sky130_fd_sc_hd__a22o_1
X_2112_ _2088_/X _2110_/Y _2111_/X _2099_/X _2747_/Q vssd1 vssd1 vccd1 vccd1 _2747_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2043_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2043_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1827_ _2052_/B _1829_/B _1887_/A vssd1 vssd1 vccd1 vccd1 _1834_/B sky130_fd_sc_hd__o21a_1
X_1689_ _1711_/A _1711_/B vssd1 vssd1 vccd1 vccd1 _1739_/A sky130_fd_sc_hd__xnor2_2
X_1758_ _1758_/A _1758_/B vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__and2_2
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2661_ _2673_/CLK _2661_/D vssd1 vssd1 vccd1 vccd1 _2661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2730_ _2769_/CLK _2730_/D _2447_/Y vssd1 vssd1 vccd1 vccd1 _2730_/Q sky130_fd_sc_hd__dfrtp_1
X_1612_ _1612_/A _1612_/B vssd1 vssd1 vccd1 vccd1 _1612_/Y sky130_fd_sc_hd__nand2_1
X_1474_ _1474_/A _1898_/B vssd1 vssd1 vccd1 vccd1 _1474_/Y sky130_fd_sc_hd__xnor2_1
X_1543_ _1687_/A vssd1 vssd1 vccd1 vccd1 _1902_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2592_ _2610_/A _2610_/B vssd1 vssd1 vccd1 vccd1 _2611_/A sky130_fd_sc_hd__nor2_1
X_2819__22 vssd1 vssd1 vccd1 vccd1 _2819__22/HI o_io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2026_ _2026_/A _2026_/B vssd1 vssd1 vccd1 vccd1 _2026_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2713_ _2757_/CLK _2713_/D vssd1 vssd1 vccd1 vccd1 _2713_/Q sky130_fd_sc_hd__dfxtp_1
X_2644_ _2601_/A _2642_/X _2643_/X _2806_/Q vssd1 vssd1 vccd1 vccd1 _2645_/B sky130_fd_sc_hd__a22o_1
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1457_ _1458_/A _1591_/A _1458_/B vssd1 vssd1 vccd1 vccd1 _1457_/Y sky130_fd_sc_hd__a21oi_1
X_1526_ _1544_/A vssd1 vssd1 vccd1 vccd1 _1901_/B sky130_fd_sc_hd__clkbuf_2
X_2575_ _2575_/A vssd1 vssd1 vccd1 vccd1 _2797_/D sky130_fd_sc_hd__clkbuf_1
X_1388_ _2065_/A _1388_/B vssd1 vssd1 vccd1 vccd1 _1388_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2009_ _2003_/A _2006_/Y _2007_/X _2008_/X vssd1 vssd1 vccd1 vccd1 _2768_/D sky130_fd_sc_hd__o31a_1
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2291_ _2669_/Q _2293_/C vssd1 vssd1 vccd1 vccd1 _2669_/D sky130_fd_sc_hd__xor2_1
X_2360_ _2503_/A vssd1 vssd1 vccd1 vccd1 _2444_/A sky130_fd_sc_hd__buf_2
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2627_ _2801_/Q _2249_/A _2625_/X _2626_/X vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__a211o_1
X_1509_ _2742_/Q vssd1 vssd1 vccd1 vccd1 _2057_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2558_ _2775_/Q vssd1 vssd1 vccd1 vccd1 _2598_/A sky130_fd_sc_hd__buf_2
X_2489_ _2489_/A vssd1 vssd1 vccd1 vccd1 _2494_/A sky130_fd_sc_hd__buf_2
XFILLER_55_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _1857_/A _1948_/A _1849_/B vssd1 vssd1 vccd1 vccd1 _1860_/Y sky130_fd_sc_hd__a21oi_1
X_1791_ _1767_/X _1791_/B _1791_/C vssd1 vssd1 vccd1 vccd1 _1791_/X sky130_fd_sc_hd__and3b_1
X_2343_ _2690_/Q _2343_/B vssd1 vssd1 vccd1 vccd1 _2343_/Y sky130_fd_sc_hd__nor2_1
X_2274_ _2274_/A vssd1 vssd1 vccd1 vccd1 _2663_/D sky130_fd_sc_hd__clkbuf_1
X_2412_ _2414_/C _2412_/B vssd1 vssd1 vccd1 vccd1 _2714_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1989_ _1992_/B _2031_/A vssd1 vssd1 vccd1 vccd1 _1989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1912_ _1912_/A _1914_/A vssd1 vssd1 vccd1 vccd1 _1913_/B sky130_fd_sc_hd__and2_1
X_1843_ _1851_/A _1852_/A vssd1 vssd1 vccd1 vccd1 _1854_/A sky130_fd_sc_hd__nand2_1
X_1774_ _1786_/A _2001_/A vssd1 vssd1 vccd1 vccd1 _1775_/B sky130_fd_sc_hd__nand2_2
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2257_ _2277_/D vssd1 vssd1 vccd1 vccd1 _2262_/A sky130_fd_sc_hd__clkbuf_2
X_2326_ _2326_/A _2328_/B vssd1 vssd1 vccd1 vccd1 _2683_/D sky130_fd_sc_hd__nor2_1
X_2188_ _2511_/A _2188_/B vssd1 vssd1 vccd1 vccd1 _2777_/D sky130_fd_sc_hd__nor2_1
XFILLER_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1490_ _1490_/A _1490_/B vssd1 vssd1 vccd1 vccd1 _1490_/Y sky130_fd_sc_hd__xnor2_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2111_ _2115_/A _2117_/A _2747_/Q vssd1 vssd1 vccd1 vccd1 _2111_/X sky130_fd_sc_hd__a21o_1
X_2042_ _2692_/D _2068_/B _2693_/Q vssd1 vssd1 vccd1 vccd1 _2137_/A sky130_fd_sc_hd__and3b_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1826_ _2732_/Q vssd1 vssd1 vccd1 vccd1 _2052_/B sky130_fd_sc_hd__clkbuf_2
X_1688_ _1688_/A _1688_/B vssd1 vssd1 vccd1 vccd1 _1711_/B sky130_fd_sc_hd__and2_1
X_1757_ _1744_/A _1756_/X _1728_/X vssd1 vssd1 vccd1 vccd1 _1758_/B sky130_fd_sc_hd__o21ai_1
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2309_ _2676_/Q _2311_/C vssd1 vssd1 vccd1 vccd1 _2676_/D sky130_fd_sc_hd__xor2_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2660_ _2673_/CLK _2660_/D vssd1 vssd1 vccd1 vccd1 _2660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1611_ _1618_/A _1618_/B vssd1 vssd1 vccd1 vccd1 _1611_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1473_ _1473_/A vssd1 vssd1 vccd1 vccd1 _1898_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1542_ _1537_/X _1538_/Y _1541_/X vssd1 vssd1 vccd1 vccd1 _1687_/A sky130_fd_sc_hd__a21o_1
XFILLER_5_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2591_ _2590_/A _2587_/Y _2590_/X vssd1 vssd1 vccd1 vccd1 _2610_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2025_ _2025_/A _2025_/B vssd1 vssd1 vccd1 vccd1 _2026_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2789_ _2793_/CLK _2789_/D vssd1 vssd1 vccd1 vccd1 _2789_/Q sky130_fd_sc_hd__dfxtp_1
X_1809_ _1807_/A _1904_/A _1778_/A vssd1 vssd1 vccd1 vccd1 _1809_/X sky130_fd_sc_hd__a21o_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2712_ _2757_/CLK _2712_/D vssd1 vssd1 vccd1 vccd1 _2712_/Q sky130_fd_sc_hd__dfxtp_1
X_2643_ _2576_/X _2183_/Y _2625_/A vssd1 vssd1 vccd1 vccd1 _2643_/X sky130_fd_sc_hd__a21o_1
X_2574_ _2645_/A _2574_/B vssd1 vssd1 vccd1 vccd1 _2575_/A sky130_fd_sc_hd__and2_1
X_1456_ _1456_/A _1456_/B vssd1 vssd1 vccd1 vccd1 _1458_/B sky130_fd_sc_hd__nor2_1
X_1525_ _1518_/A _1520_/S _1518_/B vssd1 vssd1 vccd1 vccd1 _1544_/A sky130_fd_sc_hd__a21oi_2
X_1387_ _2755_/Q vssd1 vssd1 vccd1 vccd1 _2065_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2008_ _2170_/A _2768_/Q vssd1 vssd1 vccd1 vccd1 _2008_/X sky130_fd_sc_hd__or2_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2290_ _2668_/Q _2288_/B _2289_/Y _2482_/B vssd1 vssd1 vccd1 vccd1 _2668_/D sky130_fd_sc_hd__o211a_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2557_ _2557_/A vssd1 vssd1 vccd1 vccd1 _2793_/D sky130_fd_sc_hd__clkbuf_1
X_2626_ _2802_/Q _2629_/S _2590_/X _2582_/B _2242_/A vssd1 vssd1 vccd1 vccd1 _2626_/X
+ sky130_fd_sc_hd__o221a_1
X_1439_ _1557_/B _1557_/C vssd1 vssd1 vccd1 vccd1 _1563_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1508_ _1512_/A vssd1 vssd1 vccd1 vccd1 _1749_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2488_ _2488_/A vssd1 vssd1 vccd1 vccd1 _2488_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1790_ _1767_/B _1767_/C _1760_/B _1792_/A vssd1 vssd1 vccd1 vccd1 _1791_/C sky130_fd_sc_hd__a31o_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2411_ _2714_/Q _2411_/B vssd1 vssd1 vccd1 vccd1 _2412_/B sky130_fd_sc_hd__nor2_1
X_2342_ _2688_/Q _2689_/Q _2342_/C vssd1 vssd1 vccd1 vccd1 _2342_/Y sky130_fd_sc_hd__nand3_1
X_2273_ _2275_/B _2273_/B _2285_/A vssd1 vssd1 vccd1 vccd1 _2274_/A sky130_fd_sc_hd__and3_1
XFILLER_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1988_ _1978_/Y _1979_/X _2031_/A _1975_/Y vssd1 vssd1 vccd1 vccd1 _1988_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2609_ _2609_/A vssd1 vssd1 vccd1 vccd1 _2799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1911_ _1920_/A _1803_/A _1913_/A _1912_/A _1819_/X vssd1 vssd1 vccd1 vccd1 _1914_/A
+ sky130_fd_sc_hd__a41o_1
X_1842_ _1842_/A _1842_/B vssd1 vssd1 vccd1 vccd1 _1852_/A sky130_fd_sc_hd__xor2_1
X_1773_ _1754_/X _1755_/Y _1758_/X vssd1 vssd1 vccd1 vccd1 _1786_/A sky130_fd_sc_hd__a21oi_4
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2256_ _2662_/Q _2258_/B vssd1 vssd1 vccd1 vccd1 _2277_/D sky130_fd_sc_hd__and2_1
X_2325_ _2682_/Q _2683_/Q _2325_/C vssd1 vssd1 vccd1 vccd1 _2328_/B sky130_fd_sc_hd__and3_1
X_2187_ _2527_/A _2183_/Y _2186_/X vssd1 vssd1 vccd1 vccd1 _2188_/B sky130_fd_sc_hd__a21oi_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2110_ _2110_/A vssd1 vssd1 vccd1 vccd1 _2110_/Y sky130_fd_sc_hd__inv_2
X_2041_ _2041_/A _2041_/B vssd1 vssd1 vccd1 vccd1 _2068_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1756_ _1756_/A _1756_/B vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__and2_1
X_1825_ _2731_/Q _1825_/B vssd1 vssd1 vccd1 vccd1 _1875_/A sky130_fd_sc_hd__xnor2_4
Xclkbuf_4_7_0_i_clk clkbuf_4_7_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2759_/CLK sky130_fd_sc_hd__clkbuf_2
X_2308_ _2308_/A _2311_/C vssd1 vssd1 vccd1 vccd1 _2675_/D sky130_fd_sc_hd__nor2_1
X_1687_ _1687_/A _1710_/A vssd1 vssd1 vccd1 vccd1 _1704_/B sky130_fd_sc_hd__nor2_1
X_2239_ _2511_/A _2507_/B vssd1 vssd1 vccd1 vccd1 _2776_/D sky130_fd_sc_hd__nor2_1
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1610_ _1589_/X _1599_/X _1594_/X vssd1 vssd1 vccd1 vccd1 _1618_/B sky130_fd_sc_hd__a21o_1
X_2590_ _2590_/A _2590_/B vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__or2_1
X_1472_ _1485_/A _1485_/B _1471_/X vssd1 vssd1 vccd1 vccd1 _1479_/A sky130_fd_sc_hd__o21a_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1541_ _1684_/B _1541_/B vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__and2_1
XFILLER_5_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2024_ _2024_/A vssd1 vssd1 vccd1 vccd1 _2764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1739_ _1739_/A _1739_/B vssd1 vssd1 vccd1 vccd1 _1763_/D sky130_fd_sc_hd__xnor2_1
X_2788_ _2788_/CLK _2788_/D vssd1 vssd1 vccd1 vccd1 _2788_/Q sky130_fd_sc_hd__dfxtp_1
X_1808_ _1842_/A _1841_/A vssd1 vssd1 vccd1 vccd1 _1808_/X sky130_fd_sc_hd__and2_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2711_ _2757_/CLK _2711_/D vssd1 vssd1 vccd1 vccd1 _2711_/Q sky130_fd_sc_hd__dfxtp_1
X_1524_ _1524_/A _1524_/B vssd1 vssd1 vccd1 vccd1 _1527_/A sky130_fd_sc_hd__nor2_1
X_2642_ _2576_/A _2195_/X _2590_/B _2598_/X _2805_/Q vssd1 vssd1 vccd1 vccd1 _2642_/X
+ sky130_fd_sc_hd__a32o_1
X_2573_ _2797_/Q _2572_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2574_/B sky130_fd_sc_hd__mux2_1
X_1455_ _1445_/X _1447_/X _1450_/X vssd1 vssd1 vccd1 vccd1 _1591_/A sky130_fd_sc_hd__a21o_1
X_1386_ _1394_/B _1395_/S _1394_/A vssd1 vssd1 vccd1 vccd1 _1555_/A sky130_fd_sc_hd__a21o_2
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2007_ _2006_/B _2013_/B _2006_/D _2006_/A vssd1 vssd1 vccd1 vccd1 _2007_/X sky130_fd_sc_hd__o31a_1
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_i_clk clkbuf_3_5_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1507_ _2743_/Q vssd1 vssd1 vccd1 vccd1 _2058_/A sky130_fd_sc_hd__clkbuf_2
X_2487_ _2488_/A vssd1 vssd1 vccd1 vccd1 _2487_/Y sky130_fd_sc_hd__inv_2
X_2556_ _2569_/A _2556_/B vssd1 vssd1 vccd1 vccd1 _2557_/A sky130_fd_sc_hd__and2_1
X_2625_ _2625_/A vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1438_ _1444_/B vssd1 vssd1 vccd1 vccd1 _1571_/A sky130_fd_sc_hd__clkbuf_1
X_1369_ _2757_/Q _2756_/Q vssd1 vssd1 vccd1 vccd1 _1374_/C sky130_fd_sc_hd__or2_1
XFILLER_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2341_ _2689_/Q _2343_/B vssd1 vssd1 vccd1 vccd1 _2689_/D sky130_fd_sc_hd__xnor2_1
X_2410_ _2714_/Q _2411_/B vssd1 vssd1 vccd1 vccd1 _2414_/C sky130_fd_sc_hd__and2_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2272_ _2272_/A _2272_/B _2272_/C _2272_/D vssd1 vssd1 vccd1 vccd1 _2285_/A sky130_fd_sc_hd__or4_1
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1987_ _1892_/X _1986_/X _1977_/Y vssd1 vssd1 vccd1 vccd1 _1987_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2608_ _2645_/A _2608_/B vssd1 vssd1 vccd1 vccd1 _2609_/A sky130_fd_sc_hd__and2_1
X_2539_ _2789_/Q _2550_/S _2538_/Y _2358_/X vssd1 vssd1 vccd1 vccd1 _2789_/D sky130_fd_sc_hd__o211a_1
XFILLER_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_i_clk clkbuf_2_1_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1910_ _1910_/A _1910_/B vssd1 vssd1 vccd1 vccd1 _1936_/A sky130_fd_sc_hd__xnor2_1
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1772_ _1793_/B _1789_/A vssd1 vssd1 vccd1 vccd1 _1819_/S sky130_fd_sc_hd__xor2_1
X_1841_ _1841_/A _1841_/B vssd1 vssd1 vccd1 vccd1 _1854_/B sky130_fd_sc_hd__xnor2_1
X_2324_ _2682_/Q _2325_/C _2683_/Q vssd1 vssd1 vccd1 vccd1 _2326_/A sky130_fd_sc_hd__a21oi_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2255_ _2255_/A _2258_/B vssd1 vssd1 vccd1 vccd1 _2661_/D sky130_fd_sc_hd__nor2_1
X_2186_ _2238_/B _2238_/C _2774_/Q vssd1 vssd1 vccd1 vccd1 _2186_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_4_3_0_i_clk clkbuf_4_3_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2809_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2040_ _2132_/A _2039_/X _1375_/C _1360_/B _1339_/C vssd1 vssd1 vccd1 vccd1 _2041_/B
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1686_ _1902_/A _1688_/B vssd1 vssd1 vccd1 vccd1 _1710_/A sky130_fd_sc_hd__xor2_1
X_1824_ _2730_/Q _1887_/B _1887_/A vssd1 vssd1 vccd1 vccd1 _1825_/B sky130_fd_sc_hd__o21a_1
X_1755_ _1756_/A _1755_/B vssd1 vssd1 vccd1 vccd1 _1755_/Y sky130_fd_sc_hd__xnor2_2
X_2307_ _2674_/Q _2673_/Q _2675_/Q _2307_/D vssd1 vssd1 vccd1 vccd1 _2311_/C sky130_fd_sc_hd__and4_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2238_ _2238_/A _2238_/B _2238_/C vssd1 vssd1 vccd1 vccd1 _2507_/B sky130_fd_sc_hd__or3_1
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2169_ _2693_/Q _2068_/B _2694_/Q vssd1 vssd1 vccd1 vccd1 _2693_/D sky130_fd_sc_hd__a21o_1
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1540_ _1684_/A _1539_/X _1529_/X vssd1 vssd1 vccd1 vccd1 _1541_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1471_ _1471_/A _1471_/B vssd1 vssd1 vccd1 vccd1 _1471_/X sky130_fd_sc_hd__and2_1
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2023_ _2764_/Q _2022_/Y _2032_/S vssd1 vssd1 vccd1 vccd1 _2024_/A sky130_fd_sc_hd__mux2_1
X_1807_ _1807_/A _1807_/B vssd1 vssd1 vccd1 vccd1 _1841_/A sky130_fd_sc_hd__xor2_1
X_1669_ _1669_/A _1669_/B vssd1 vssd1 vccd1 vccd1 _1669_/X sky130_fd_sc_hd__xor2_1
X_1738_ _1767_/A _1764_/B _1731_/B _1737_/Y vssd1 vssd1 vccd1 vccd1 _1739_/B sky130_fd_sc_hd__a31o_1
X_2787_ _2788_/CLK _2787_/D vssd1 vssd1 vccd1 vccd1 _2787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_0_0_i_clk clkbuf_3_1_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2710_ _2757_/CLK _2710_/D vssd1 vssd1 vccd1 vccd1 _2710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1454_ _2104_/A _1454_/B vssd1 vssd1 vccd1 vccd1 _1461_/A sky130_fd_sc_hd__xnor2_1
X_1523_ _1539_/A vssd1 vssd1 vccd1 vccd1 _1523_/Y sky130_fd_sc_hd__inv_2
X_2641_ _2805_/Q _2617_/X _2640_/X _2636_/X vssd1 vssd1 vccd1 vccd1 _2805_/D sky130_fd_sc_hd__o211a_1
X_2572_ _2769_/Q _2796_/Q _2598_/A vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__mux2_1
X_1385_ _1390_/A _1549_/A vssd1 vssd1 vccd1 vccd1 _1394_/A sky130_fd_sc_hd__and2b_1
XFILLER_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2006_ _2006_/A _2006_/B _2013_/B _2006_/D vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__nor4_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2624_ _2801_/Q _2617_/X _2623_/X _2358_/X vssd1 vssd1 vccd1 vccd1 _2801_/D sky130_fd_sc_hd__o211a_1
X_1437_ _1446_/A _1446_/B _1444_/A _1448_/A _1448_/B vssd1 vssd1 vccd1 vccd1 _1444_/B
+ sky130_fd_sc_hd__o311ai_1
X_1506_ _1506_/A _1545_/A _1545_/B vssd1 vssd1 vccd1 vccd1 _1524_/B sky130_fd_sc_hd__and3_1
X_2486_ _2488_/A vssd1 vssd1 vccd1 vccd1 _2486_/Y sky130_fd_sc_hd__inv_2
X_2555_ _2793_/Q _2553_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2556_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1368_ _2758_/Q vssd1 vssd1 vccd1 vccd1 _2075_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _2340_/A vssd1 vssd1 vccd1 vccd1 _2688_/D sky130_fd_sc_hd__clkbuf_1
X_2271_ _2271_/A _2271_/B _2271_/C _2271_/D vssd1 vssd1 vccd1 vccd1 _2272_/D sky130_fd_sc_hd__or4_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ _1991_/A _1992_/A _1992_/B _1983_/X _1985_/A vssd1 vssd1 vccd1 vccd1 _1986_/X
+ sky130_fd_sc_hd__a311o_1
X_2607_ _2799_/Q _2597_/X _2606_/X _2601_/A vssd1 vssd1 vccd1 vccd1 _2608_/B sky130_fd_sc_hd__a22o_1
X_2469_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2469_/Y sky130_fd_sc_hd__inv_2
X_2538_ _2537_/Y _2249_/A _2550_/S vssd1 vssd1 vccd1 vccd1 _2538_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1840_ _1842_/A _1842_/B vssd1 vssd1 vccd1 vccd1 _1841_/B sky130_fd_sc_hd__nand2_1
X_1771_ _1793_/A _1793_/C _2001_/A vssd1 vssd1 vccd1 vccd1 _1789_/A sky130_fd_sc_hd__and3_1
X_2254_ _2660_/Q _2659_/Q _2661_/Q vssd1 vssd1 vccd1 vccd1 _2258_/B sky130_fd_sc_hd__and3_1
X_2323_ _2682_/Q _2325_/C vssd1 vssd1 vccd1 vccd1 _2682_/D sky130_fd_sc_hd__xor2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2185_ _2785_/Q _2784_/Q _2783_/Q _2782_/Q vssd1 vssd1 vccd1 vccd1 _2238_/C sky130_fd_sc_hd__or4_1
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1969_ _1977_/B vssd1 vssd1 vccd1 vccd1 _1978_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1823_ _1823_/A vssd1 vssd1 vccd1 vccd1 _1887_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1685_ _1685_/A _1685_/B vssd1 vssd1 vccd1 vccd1 _1704_/A sky130_fd_sc_hd__xnor2_1
X_1754_ _1744_/A _1746_/Y _1728_/X _1755_/B _1753_/Y vssd1 vssd1 vccd1 vccd1 _1754_/X
+ sky130_fd_sc_hd__a311o_2
X_2306_ _2674_/Q _2304_/B _2675_/Q vssd1 vssd1 vccd1 vccd1 _2308_/A sky130_fd_sc_hd__a21oi_1
X_2237_ _2774_/Q vssd1 vssd1 vccd1 vccd1 _2238_/A sky130_fd_sc_hd__clkinv_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2099_ _2099_/A vssd1 vssd1 vccd1 vccd1 _2099_/X sky130_fd_sc_hd__clkbuf_2
X_2168_ _2168_/A vssd1 vssd1 vccd1 vccd1 _2728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1470_ _1470_/A _1470_/B _1470_/C vssd1 vssd1 vccd1 vccd1 _1471_/B sky130_fd_sc_hd__or3_1
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2022_ _2022_/A _2022_/B vssd1 vssd1 vccd1 vccd1 _2022_/Y sky130_fd_sc_hd__xnor2_1
X_2786_ _2788_/CLK _2786_/D vssd1 vssd1 vccd1 vccd1 _2786_/Q sky130_fd_sc_hd__dfxtp_1
X_1806_ _2054_/A _1806_/B vssd1 vssd1 vccd1 vccd1 _1842_/A sky130_fd_sc_hd__xor2_2
X_1599_ _1599_/A _1613_/B vssd1 vssd1 vccd1 vccd1 _1599_/X sky130_fd_sc_hd__or2b_1
X_1668_ _1655_/A _1667_/A _1655_/B vssd1 vssd1 vccd1 vccd1 _1669_/B sky130_fd_sc_hd__o21ba_1
X_1737_ _1737_/A vssd1 vssd1 vccd1 vccd1 _1737_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2640_ _2804_/Q _2248_/A _2639_/X _2244_/A _2625_/X vssd1 vssd1 vccd1 vccd1 _2640_/X
+ sky130_fd_sc_hd__a221o_1
X_1453_ _2748_/Q vssd1 vssd1 vccd1 vccd1 _2104_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1522_ _2057_/A _1522_/B vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__xor2_1
X_2571_ _2571_/A vssd1 vssd1 vccd1 vccd1 _2645_/A sky130_fd_sc_hd__clkbuf_2
X_1384_ _1365_/Y _1383_/B _1549_/B vssd1 vssd1 vccd1 vccd1 _1395_/S sky130_fd_sc_hd__o21ai_1
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2005_ _2030_/A _2005_/B vssd1 vssd1 vccd1 vccd1 _2006_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2769_ _2769_/CLK _2769_/D _2493_/Y vssd1 vssd1 vccd1 vccd1 _2769_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2554_ _2554_/A vssd1 vssd1 vccd1 vccd1 _2573_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2623_ _2625_/A _2623_/B _2622_/X vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__or3b_1
X_1436_ _1440_/A _1557_/B _1433_/Y vssd1 vssd1 vccd1 vccd1 _1448_/B sky130_fd_sc_hd__o21ai_1
X_1367_ _2756_/Q _1376_/B vssd1 vssd1 vccd1 vccd1 _1367_/Y sky130_fd_sc_hd__xnor2_1
X_1505_ _1545_/A _1545_/B _1506_/A vssd1 vssd1 vccd1 vccd1 _1524_/A sky130_fd_sc_hd__a21oi_1
X_2485_ _2488_/A vssd1 vssd1 vccd1 vccd1 _2485_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2270_ _2664_/Q _2663_/Q _2270_/C _2269_/X vssd1 vssd1 vccd1 vccd1 _2271_/D sky130_fd_sc_hd__or4b_1
X_1985_ _1985_/A _2031_/A vssd1 vssd1 vccd1 vccd1 _1985_/X sky130_fd_sc_hd__and2_1
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2606_ _2576_/A _2580_/Y _2605_/Y _2598_/X _2798_/Q vssd1 vssd1 vccd1 vccd1 _2606_/X
+ sky130_fd_sc_hd__a32o_1
X_2537_ _2761_/Q vssd1 vssd1 vccd1 vccd1 _2537_/Y sky130_fd_sc_hd__inv_2
X_1419_ _2751_/Q _1419_/B vssd1 vssd1 vccd1 vccd1 _1428_/A sky130_fd_sc_hd__xor2_2
X_2468_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2468_/Y sky130_fd_sc_hd__inv_2
X_2399_ _2709_/Q _2400_/C vssd1 vssd1 vccd1 vccd1 _2709_/D sky130_fd_sc_hd__xor2_1
XFILLER_22_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1770_ _1793_/D vssd1 vssd1 vccd1 vccd1 _2001_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2253_ _2660_/Q _2659_/Q _2661_/Q vssd1 vssd1 vccd1 vccd1 _2255_/A sky130_fd_sc_hd__a21oi_1
X_2322_ _2322_/A _2325_/C vssd1 vssd1 vccd1 vccd1 _2681_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2184_ _2780_/Q _2779_/Q _2778_/Q _2781_/Q vssd1 vssd1 vccd1 vccd1 _2238_/B sky130_fd_sc_hd__or4b_1
X_1899_ _1899_/A _1899_/B _1899_/C _1898_/X vssd1 vssd1 vccd1 vccd1 _1900_/B sky130_fd_sc_hd__or4b_1
X_1968_ _1983_/A _1971_/A _1991_/A _1971_/B _1967_/Y vssd1 vssd1 vccd1 vccd1 _1977_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1822_ _1894_/A _2728_/Q vssd1 vssd1 vccd1 vccd1 _1887_/B sky130_fd_sc_hd__or2_1
XFILLER_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1753_ _1776_/A vssd1 vssd1 vccd1 vccd1 _1753_/Y sky130_fd_sc_hd__inv_2
X_1684_ _1684_/A _1684_/B _1688_/B vssd1 vssd1 vccd1 vccd1 _1685_/B sky130_fd_sc_hd__and3_1
X_2305_ _2674_/Q _2304_/B _2304_/Y _2482_/B vssd1 vssd1 vccd1 vccd1 _2674_/D sky130_fd_sc_hd__o211a_1
X_2236_ _2236_/A vssd1 vssd1 vccd1 vccd1 _2658_/D sky130_fd_sc_hd__clkbuf_1
X_2167_ _2113_/A _2099_/A _2728_/Q vssd1 vssd1 vccd1 vccd1 _2168_/A sky130_fd_sc_hd__mux2_1
X_2098_ _2102_/A _2102_/B _2751_/Q vssd1 vssd1 vccd1 vccd1 _2098_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2021_ _2026_/A _2025_/B _2025_/A vssd1 vssd1 vccd1 vccd1 _2022_/B sky130_fd_sc_hd__o21ai_1
XFILLER_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1736_ _1764_/B _1764_/C _1735_/Y vssd1 vssd1 vccd1 vccd1 _1762_/A sky130_fd_sc_hd__a21oi_1
X_2785_ _2793_/CLK _2785_/D vssd1 vssd1 vccd1 vccd1 _2785_/Q sky130_fd_sc_hd__dfxtp_1
X_1805_ _1823_/A _1805_/B vssd1 vssd1 vccd1 vccd1 _1806_/B sky130_fd_sc_hd__nand2_1
X_1598_ _1620_/A _1619_/A _1619_/B _1591_/B _1597_/X vssd1 vssd1 vccd1 vccd1 _1613_/B
+ sky130_fd_sc_hd__a41o_1
X_1667_ _1667_/A _1667_/B vssd1 vssd1 vccd1 vccd1 _1691_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2219_ _2219_/A _2233_/C vssd1 vssd1 vccd1 vccd1 _2228_/A sky130_fd_sc_hd__nand2_2
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2816__19 vssd1 vssd1 vccd1 vccd1 _2816__19/HI o_io_oeb[5] sky130_fd_sc_hd__conb_1
X_2570_ _2570_/A vssd1 vssd1 vccd1 vccd1 _2796_/D sky130_fd_sc_hd__clkbuf_1
X_1452_ _1458_/A _1473_/A vssd1 vssd1 vccd1 vccd1 _1462_/A sky130_fd_sc_hd__xnor2_1
X_1383_ _1392_/A _1383_/B _1383_/C vssd1 vssd1 vccd1 vccd1 _1394_/B sky130_fd_sc_hd__or3_1
X_1521_ _1677_/A vssd1 vssd1 vccd1 vccd1 _1684_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2004_ _2170_/A _1998_/X _2001_/X _2003_/X vssd1 vssd1 vccd1 vccd1 _2769_/D sky130_fd_sc_hd__a31o_1
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2699_ _2806_/CLK _2699_/D vssd1 vssd1 vccd1 vccd1 _2699_/Q sky130_fd_sc_hd__dfxtp_1
X_1719_ _1719_/A _1719_/B vssd1 vssd1 vccd1 vccd1 _1767_/B sky130_fd_sc_hd__xor2_2
X_2768_ _2769_/CLK _2768_/D _2492_/Y vssd1 vssd1 vccd1 vccd1 _2768_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1504_ _1504_/A vssd1 vssd1 vccd1 vccd1 _1506_/A sky130_fd_sc_hd__inv_2
X_2553_ _2765_/Q _2792_/Q _2553_/S vssd1 vssd1 vccd1 vccd1 _2553_/X sky130_fd_sc_hd__mux2_1
X_2622_ _2622_/A _2638_/A _2622_/C _2576_/X vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__or4b_1
X_1435_ _1435_/A vssd1 vssd1 vccd1 vccd1 _1557_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1366_ _1341_/B _1360_/B _1374_/B _1373_/A vssd1 vssd1 vccd1 vccd1 _1376_/B sky130_fd_sc_hd__o31a_1
X_2484_ _2488_/A vssd1 vssd1 vccd1 vccd1 _2484_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1984_ _1991_/A _1992_/A _1992_/B _1983_/X vssd1 vssd1 vccd1 vccd1 _2031_/A sky130_fd_sc_hd__a31o_1
X_2467_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2467_/Y sky130_fd_sc_hd__inv_2
X_2536_ _2554_/A vssd1 vssd1 vccd1 vccd1 _2550_/S sky130_fd_sc_hd__clkbuf_2
X_2605_ _2587_/Y _2590_/X _2610_/B vssd1 vssd1 vccd1 vccd1 _2605_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_57_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1349_ _1349_/A vssd1 vssd1 vccd1 vccd1 _1483_/A sky130_fd_sc_hd__inv_2
X_1418_ _1334_/A _2750_/Q _1432_/B vssd1 vssd1 vccd1 vccd1 _1419_/B sky130_fd_sc_hd__a21o_1
X_2398_ _2400_/C _2398_/B vssd1 vssd1 vccd1 vccd1 _2708_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2321_ _2681_/Q _2321_/B vssd1 vssd1 vccd1 vccd1 _2325_/C sky130_fd_sc_hd__and2_1
XFILLER_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2252_ _2660_/Q _2659_/Q vssd1 vssd1 vccd1 vccd1 _2660_/D sky130_fd_sc_hd__xor2_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2183_ _2183_/A _2183_/B vssd1 vssd1 vccd1 vccd1 _2183_/Y sky130_fd_sc_hd__nand2_2
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1898_ _1898_/A _1898_/B _1898_/C vssd1 vssd1 vccd1 vccd1 _1898_/X sky130_fd_sc_hd__and3_1
X_1967_ _1943_/X _1965_/X _1966_/Y vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__a21oi_1
X_2519_ _2519_/A _2519_/B vssd1 vssd1 vccd1 vccd1 _2785_/D sky130_fd_sc_hd__nor2_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1683_ _1691_/A _1688_/A _1711_/A _1675_/A _1682_/X vssd1 vssd1 vccd1 vccd1 _1688_/B
+ sky130_fd_sc_hd__a41o_1
X_1752_ _2055_/A _1752_/B vssd1 vssd1 vccd1 vccd1 _1776_/A sky130_fd_sc_hd__xnor2_2
X_1821_ _2729_/Q vssd1 vssd1 vccd1 vccd1 _1894_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2304_ _2674_/Q _2304_/B vssd1 vssd1 vccd1 vccd1 _2304_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2097_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2097_/Y sky130_fd_sc_hd__inv_2
X_2235_ _2235_/A _2235_/B vssd1 vssd1 vccd1 vccd1 _2236_/A sky130_fd_sc_hd__or2_1
X_2166_ _1887_/B _2165_/Y _2073_/X _2099_/A _1894_/A vssd1 vssd1 vccd1 vccd1 _2729_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2020_ _2020_/A vssd1 vssd1 vccd1 vccd1 _2765_/D sky130_fd_sc_hd__clkbuf_1
X_1666_ _1665_/Y _1661_/C _1650_/Y vssd1 vssd1 vccd1 vccd1 _1667_/B sky130_fd_sc_hd__a21boi_1
X_1735_ _1734_/A _1764_/C _1734_/B vssd1 vssd1 vccd1 vccd1 _1735_/Y sky130_fd_sc_hd__a21oi_1
X_1804_ _2736_/Q vssd1 vssd1 vccd1 vccd1 _2054_/A sky130_fd_sc_hd__clkbuf_2
X_2784_ _2793_/CLK _2784_/D vssd1 vssd1 vccd1 vccd1 _2784_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _1577_/X _1597_/B vssd1 vssd1 vccd1 vccd1 _1597_/X sky130_fd_sc_hd__and2b_1
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2218_ _2227_/A _2225_/B _2218_/C vssd1 vssd1 vccd1 vccd1 _2233_/C sky130_fd_sc_hd__or3_2
X_2149_ _2149_/A _2149_/B vssd1 vssd1 vccd1 vccd1 _2149_/X sky130_fd_sc_hd__or2_1
XFILLER_14_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1520_ _1518_/Y _1518_/A _1520_/S vssd1 vssd1 vccd1 vccd1 _1677_/A sky130_fd_sc_hd__mux2_1
X_1451_ _1445_/X _1447_/X _1450_/X vssd1 vssd1 vccd1 vccd1 _1473_/A sky130_fd_sc_hd__a21oi_1
X_1382_ _2755_/Q _1388_/B vssd1 vssd1 vccd1 vccd1 _1392_/A sky130_fd_sc_hd__xor2_2
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2003_ _2003_/A _2769_/Q vssd1 vssd1 vccd1 vccd1 _2003_/X sky130_fd_sc_hd__and2_1
X_1649_ _1900_/A _1651_/B _1635_/B vssd1 vssd1 vccd1 vccd1 _1649_/X sky130_fd_sc_hd__o21a_1
X_2698_ _2806_/CLK _2698_/D vssd1 vssd1 vccd1 vccd1 _2698_/Q sky130_fd_sc_hd__dfxtp_1
X_1718_ _1731_/A _1764_/C vssd1 vssd1 vccd1 vccd1 _1719_/B sky130_fd_sc_hd__nand2_1
X_2767_ _2769_/CLK _2767_/D _2491_/Y vssd1 vssd1 vccd1 vccd1 _2767_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1503_ _1490_/Y _1900_/A _1502_/X vssd1 vssd1 vccd1 vccd1 _1545_/B sky130_fd_sc_hd__o21a_1
X_2552_ _2552_/A vssd1 vssd1 vccd1 vccd1 _2792_/D sky130_fd_sc_hd__clkbuf_1
X_2483_ _2489_/A vssd1 vssd1 vccd1 vccd1 _2488_/A sky130_fd_sc_hd__buf_2
X_2621_ _2621_/A _2621_/B vssd1 vssd1 vccd1 vccd1 _2638_/A sky130_fd_sc_hd__or2_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1434_ _1435_/A _1431_/C _1433_/Y _1440_/A vssd1 vssd1 vccd1 vccd1 _1448_/A sky130_fd_sc_hd__a211o_1
X_1365_ _2757_/Q _1365_/B vssd1 vssd1 vccd1 vccd1 _1365_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2604_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2798_/D sky130_fd_sc_hd__clkbuf_1
X_1983_ _1983_/A _1983_/B vssd1 vssd1 vccd1 vccd1 _1983_/X sky130_fd_sc_hd__xor2_1
XFILLER_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1417_ _1334_/A _1359_/D _1454_/B vssd1 vssd1 vccd1 vccd1 _1432_/B sky130_fd_sc_hd__a21o_1
X_2466_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2466_/Y sky130_fd_sc_hd__inv_2
X_2535_ _2772_/Q _2775_/Q _2190_/X vssd1 vssd1 vccd1 vccd1 _2554_/A sky130_fd_sc_hd__o21a_1
X_1348_ _2746_/Q _1348_/B vssd1 vssd1 vccd1 vccd1 _1349_/A sky130_fd_sc_hd__xor2_2
XFILLER_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2397_ _2708_/Q _2397_/B vssd1 vssd1 vccd1 vccd1 _2398_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2251_ _2659_/Q vssd1 vssd1 vccd1 vccd1 _2659_/D sky130_fd_sc_hd__clkinv_2
X_2320_ _2681_/Q _2321_/B vssd1 vssd1 vccd1 vccd1 _2322_/A sky130_fd_sc_hd__nor2_1
X_2182_ _2632_/A _2622_/A vssd1 vssd1 vccd1 vccd1 _2183_/B sky130_fd_sc_hd__and2_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1966_ _1965_/X _2022_/A _1943_/X vssd1 vssd1 vccd1 vccd1 _1966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1897_ _1581_/A _1579_/B _1897_/C _1897_/D vssd1 vssd1 vccd1 vccd1 _1898_/C sky130_fd_sc_hd__and4bb_1
X_2518_ _2785_/Q _2784_/Q _2514_/A _2489_/A vssd1 vssd1 vccd1 vccd1 _2519_/B sky130_fd_sc_hd__a31o_1
X_2449_ _2451_/A vssd1 vssd1 vccd1 vccd1 _2449_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1820_ _1920_/A _1803_/X _1912_/A _1819_/X vssd1 vssd1 vccd1 vccd1 _2005_/B sky130_fd_sc_hd__a31oi_4
XFILLER_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1682_ _1682_/A _1682_/B vssd1 vssd1 vccd1 vccd1 _1682_/X sky130_fd_sc_hd__xor2_1
X_1751_ _1823_/A _2055_/B _1777_/B vssd1 vssd1 vccd1 vccd1 _1752_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2303_ _2673_/Q _2307_/D _2302_/Y _2482_/B vssd1 vssd1 vccd1 vccd1 _2673_/D sky130_fd_sc_hd__o211a_1
X_2234_ _2657_/D _2234_/B vssd1 vssd1 vccd1 vccd1 _2234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2096_ _2093_/B _2095_/Y _2063_/A _2086_/X vssd1 vssd1 vccd1 vccd1 _2752_/D sky130_fd_sc_hd__a2bb2o_1
X_2165_ _2165_/A vssd1 vssd1 vccd1 vccd1 _2165_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1949_ _1948_/A _2018_/A _1948_/B vssd1 vssd1 vccd1 vccd1 _1949_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2783_ _2783_/CLK _2783_/D vssd1 vssd1 vccd1 vccd1 _2783_/Q sky130_fd_sc_hd__dfxtp_1
X_1803_ _1803_/A _1913_/A vssd1 vssd1 vccd1 vccd1 _1803_/X sky130_fd_sc_hd__and2_1
X_1596_ _1576_/A _1581_/B _1577_/C _1595_/A vssd1 vssd1 vccd1 vccd1 _1597_/B sky130_fd_sc_hd__a31o_1
X_1665_ _1665_/A vssd1 vssd1 vccd1 vccd1 _1665_/Y sky130_fd_sc_hd__inv_2
X_1734_ _1734_/A _1734_/B vssd1 vssd1 vccd1 vccd1 _1764_/B sky130_fd_sc_hd__and2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2217_ _2227_/B _2221_/A vssd1 vssd1 vccd1 vccd1 _2218_/C sky130_fd_sc_hd__nand2_1
X_2079_ _2079_/A vssd1 vssd1 vccd1 vccd1 _2079_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2148_ _2149_/A _2149_/B vssd1 vssd1 vccd1 vccd1 _2148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1450_ _1448_/X _1449_/X _1571_/A vssd1 vssd1 vccd1 vccd1 _1450_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1381_ _1410_/A _2064_/A _1393_/B vssd1 vssd1 vccd1 vccd1 _1388_/B sky130_fd_sc_hd__a21o_1
X_2002_ _2695_/Q vssd1 vssd1 vccd1 vccd1 _2003_/A sky130_fd_sc_hd__inv_2
X_2766_ _2769_/CLK _2766_/D _2490_/Y vssd1 vssd1 vccd1 vccd1 _2766_/Q sky130_fd_sc_hd__dfrtp_1
X_1579_ _1559_/B _1579_/B vssd1 vssd1 vccd1 vccd1 _1579_/X sky130_fd_sc_hd__and2b_1
X_1648_ _1643_/Y _1636_/A _1647_/X _1640_/X vssd1 vssd1 vccd1 vccd1 _1651_/B sky130_fd_sc_hd__a31oi_2
X_2697_ _2807_/CLK _2697_/D vssd1 vssd1 vccd1 vccd1 _2697_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1717_ _1731_/B vssd1 vssd1 vccd1 vccd1 _1764_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2821__24 vssd1 vssd1 vccd1 vccd1 _2821__24/HI o_io_oeb[10] sky130_fd_sc_hd__conb_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2620_ _2577_/A _2611_/A _2593_/A vssd1 vssd1 vccd1 vccd1 _2621_/B sky130_fd_sc_hd__o21a_1
X_1433_ _1433_/A _1433_/B vssd1 vssd1 vccd1 vccd1 _1433_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1502_ _1490_/A _1488_/X _1492_/X vssd1 vssd1 vccd1 vccd1 _1502_/X sky130_fd_sc_hd__a21o_1
X_2482_ _2760_/Q _2482_/B vssd1 vssd1 vccd1 vccd1 _2760_/D sky130_fd_sc_hd__xnor2_1
X_2551_ _2569_/A _2551_/B vssd1 vssd1 vccd1 vccd1 _2552_/A sky130_fd_sc_hd__and2_1
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1364_ _2756_/Q _1360_/A _1360_/B _1374_/B _2759_/Q vssd1 vssd1 vccd1 vccd1 _1365_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2749_ _2758_/CLK _2749_/D _2469_/Y vssd1 vssd1 vccd1 vccd1 _2749_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1982_ _1991_/A _1972_/A _1978_/C _1981_/Y vssd1 vssd1 vccd1 vccd1 _1983_/B sky130_fd_sc_hd__a31o_1
X_2603_ _2645_/A _2603_/B vssd1 vssd1 vccd1 vccd1 _2604_/A sky130_fd_sc_hd__and2_1
X_2534_ _2534_/A vssd1 vssd1 vccd1 vccd1 _2788_/D sky130_fd_sc_hd__clkbuf_1
X_1416_ _1405_/X _1414_/X _1551_/A vssd1 vssd1 vccd1 vccd1 _1435_/A sky130_fd_sc_hd__a21bo_1
X_1347_ _2059_/A _2744_/Q _1341_/B _1334_/A vssd1 vssd1 vccd1 vccd1 _1348_/B sky130_fd_sc_hd__o31ai_2
X_2465_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2465_/Y sky130_fd_sc_hd__inv_2
X_2396_ _2708_/Q _2397_/B vssd1 vssd1 vccd1 vccd1 _2400_/C sky130_fd_sc_hd__and2_1
XFILLER_3_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2250_ _2250_/A vssd1 vssd1 vccd1 vccd1 _2774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2181_ _2581_/A vssd1 vssd1 vccd1 vccd1 _2622_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1965_ _1983_/A _1965_/B _1965_/C vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__and3_1
X_1896_ _1875_/A _1895_/X _1578_/A _1555_/Y vssd1 vssd1 vccd1 vccd1 _1897_/D sky130_fd_sc_hd__o211a_1
X_2517_ _2784_/Q _2514_/A _2785_/Q vssd1 vssd1 vccd1 vccd1 _2519_/A sky130_fd_sc_hd__a21oi_1
X_2379_ _2701_/Q _2382_/C vssd1 vssd1 vccd1 vccd1 _2380_/C sky130_fd_sc_hd__or2_1
X_2448_ _2451_/A vssd1 vssd1 vccd1 vccd1 _2448_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1750_ _2736_/Q _1805_/B _1823_/A vssd1 vssd1 vccd1 vccd1 _1777_/B sky130_fd_sc_hd__o21a_1
X_1681_ _1671_/A _1691_/A _1679_/B _1667_/A vssd1 vssd1 vccd1 vccd1 _1682_/B sky130_fd_sc_hd__a31o_1
X_2302_ _2304_/B vssd1 vssd1 vccd1 vccd1 _2302_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2233_ _2230_/X _2233_/B _2233_/C vssd1 vssd1 vccd1 vccd1 _2233_/Y sky130_fd_sc_hd__nand3b_4
X_2164_ _2043_/X _2162_/Y _2163_/X _2146_/X _2163_/A vssd1 vssd1 vccd1 vccd1 _2730_/D
+ sky130_fd_sc_hd__a32o_1
X_2095_ _2063_/A _2097_/A _2043_/X vssd1 vssd1 vccd1 vccd1 _2095_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1948_ _1948_/A _1948_/B vssd1 vssd1 vccd1 vccd1 _1948_/Y sky130_fd_sc_hd__nor2_1
X_1879_ _1879_/A _1879_/B vssd1 vssd1 vccd1 vccd1 _1883_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1733_ _1733_/A vssd1 vssd1 vccd1 vccd1 _1767_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2782_ _2783_/CLK _2782_/D vssd1 vssd1 vccd1 vccd1 _2782_/Q sky130_fd_sc_hd__dfxtp_1
X_1802_ _1802_/A _1802_/B vssd1 vssd1 vccd1 vccd1 _1913_/A sky130_fd_sc_hd__xnor2_2
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ _1595_/A _1620_/A _1619_/A _1619_/B vssd1 vssd1 vccd1 vccd1 _1599_/A sky130_fd_sc_hd__and4_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1664_ _1656_/Y _1658_/X _1650_/Y _1665_/A vssd1 vssd1 vccd1 vccd1 _1667_/A sky130_fd_sc_hd__a211oi_2
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2216_ _2216_/A vssd1 vssd1 vccd1 vccd1 _2225_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2147_ _2137_/X _2144_/Y _2145_/X _2146_/X _2054_/A vssd1 vssd1 vccd1 vccd1 _2736_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2078_ _2073_/X _2074_/Y _2075_/X _2077_/X _2075_/A vssd1 vssd1 vccd1 vccd1 _2758_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1380_ _2753_/Q _2752_/Q _1410_/B _1373_/A vssd1 vssd1 vccd1 vccd1 _1393_/B sky130_fd_sc_hd__o31a_1
X_2001_ _2001_/A _2013_/B _2006_/B _1909_/X vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__or4b_1
XFILLER_50_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2696_ _2806_/CLK _2696_/D vssd1 vssd1 vccd1 vccd1 _2696_/Q sky130_fd_sc_hd__dfxtp_1
X_1716_ _1703_/Y _1733_/A _1734_/A _1734_/B _1715_/X vssd1 vssd1 vccd1 vccd1 _1731_/B
+ sky130_fd_sc_hd__a41o_1
X_2765_ _2769_/CLK _2765_/D _2488_/Y vssd1 vssd1 vccd1 vccd1 _2765_/Q sky130_fd_sc_hd__dfrtp_1
X_1578_ _1578_/A _1578_/B vssd1 vssd1 vccd1 vccd1 _1578_/X sky130_fd_sc_hd__and2_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1647_ _1658_/A _1669_/A vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__and2b_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2550_ _2792_/Q _2549_/X _2550_/S vssd1 vssd1 vccd1 vccd1 _2551_/B sky130_fd_sc_hd__mux2_1
X_1432_ _2750_/Q _1432_/B vssd1 vssd1 vccd1 vccd1 _1444_/A sky130_fd_sc_hd__xor2_2
X_1501_ _1501_/A vssd1 vssd1 vccd1 vccd1 _1900_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1363_ _2755_/Q _2754_/Q _2753_/Q _2752_/Q vssd1 vssd1 vccd1 vccd1 _1374_/B sky130_fd_sc_hd__or4_2
X_2481_ _2481_/A vssd1 vssd1 vccd1 vccd1 _2481_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2679_ _2727_/CLK _2679_/D vssd1 vssd1 vccd1 vccd1 _2679_/Q sky130_fd_sc_hd__dfxtp_1
X_2748_ _2758_/CLK _2748_/D _2468_/Y vssd1 vssd1 vccd1 vccd1 _2748_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1981_ _1981_/A vssd1 vssd1 vccd1 vccd1 _1981_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2602_ _2798_/Q _2597_/X _2599_/X _2655_/B vssd1 vssd1 vccd1 vccd1 _2603_/B sky130_fd_sc_hd__a22o_1
X_2533_ _2531_/X _2533_/B vssd1 vssd1 vccd1 vccd1 _2534_/A sky130_fd_sc_hd__and2b_1
X_1415_ _1409_/Y _1411_/X _1405_/X vssd1 vssd1 vccd1 vccd1 _1551_/A sky130_fd_sc_hd__a21o_1
X_1346_ _1488_/B vssd1 vssd1 vccd1 vccd1 _1494_/A sky130_fd_sc_hd__inv_2
X_2464_ _2470_/A vssd1 vssd1 vccd1 vccd1 _2469_/A sky130_fd_sc_hd__buf_2
X_2395_ _2397_/B _2395_/B vssd1 vssd1 vccd1 vccd1 _2707_/D sky130_fd_sc_hd__nor2_1
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2180_ _2787_/Q vssd1 vssd1 vccd1 vccd1 _2581_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1895_ _2041_/A _1893_/Y _1888_/B _2165_/A _1888_/X vssd1 vssd1 vccd1 vccd1 _1895_/X
+ sky130_fd_sc_hd__o221a_1
X_1964_ _1964_/A _1964_/B vssd1 vssd1 vccd1 vccd1 _1971_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2516_ _2784_/Q _2514_/A _2515_/Y vssd1 vssd1 vccd1 vccd1 _2784_/D sky130_fd_sc_hd__o21a_1
X_2447_ _2451_/A vssd1 vssd1 vccd1 vccd1 _2447_/Y sky130_fd_sc_hd__inv_2
X_2378_ _2383_/B vssd1 vssd1 vccd1 vccd1 _2380_/B sky130_fd_sc_hd__clkinv_2
X_1329_ _1329_/A vssd1 vssd1 vccd1 vccd1 _2694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2301_ _2673_/Q _2307_/D vssd1 vssd1 vccd1 vccd1 _2304_/B sky130_fd_sc_hd__and2_1
X_1680_ _1680_/A _1680_/B vssd1 vssd1 vccd1 vccd1 _1711_/A sky130_fd_sc_hd__xnor2_2
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2232_ _2222_/B _2225_/C _2233_/B vssd1 vssd1 vccd1 vccd1 _2232_/X sky130_fd_sc_hd__a21bo_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2163_ _2163_/A _2165_/A vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__or2_1
XFILLER_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2094_ _2088_/X _2092_/Y _2093_/X _2077_/X _2093_/A vssd1 vssd1 vccd1 vccd1 _2753_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1947_ _1947_/A _1964_/A vssd1 vssd1 vccd1 vccd1 _1965_/B sky130_fd_sc_hd__or2_1
X_1878_ _1878_/A _1878_/B vssd1 vssd1 vccd1 vccd1 _1879_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_12_0_i_clk clkbuf_3_6_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _2757_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1663_ _1672_/A _1680_/A _1661_/X _1662_/Y vssd1 vssd1 vccd1 vccd1 _1671_/A sky130_fd_sc_hd__o22a_1
X_1732_ _1903_/A _1745_/A vssd1 vssd1 vccd1 vccd1 _1767_/C sky130_fd_sc_hd__or2_1
X_2781_ _2783_/CLK _2781_/D vssd1 vssd1 vccd1 vccd1 _2781_/Q sky130_fd_sc_hd__dfxtp_1
X_1801_ _1904_/A _1801_/B vssd1 vssd1 vccd1 vccd1 _1802_/B sky130_fd_sc_hd__or2_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _1612_/A _1612_/B _1614_/A _1614_/B vssd1 vssd1 vccd1 vccd1 _1594_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2077_ _2099_/A vssd1 vssd1 vccd1 vccd1 _2077_/X sky130_fd_sc_hd__clkbuf_2
X_2215_ _2222_/A _2215_/B vssd1 vssd1 vccd1 vccd1 _2219_/A sky130_fd_sc_hd__nand2_1
X_2146_ _2146_/A vssd1 vssd1 vccd1 vccd1 _2146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2000_ _2030_/A _2013_/A vssd1 vssd1 vccd1 vccd1 _2006_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1646_ _1639_/D _1642_/B _1645_/Y vssd1 vssd1 vccd1 vccd1 _1669_/A sky130_fd_sc_hd__a21boi_1
X_1715_ _1712_/Y _1713_/X _1713_/A _1714_/X vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__o2bb2a_1
X_2764_ _2769_/CLK _2764_/D _2487_/Y vssd1 vssd1 vccd1 vccd1 _2764_/Q sky130_fd_sc_hd__dfrtp_1
X_2695_ _2805_/CLK _2695_/D _2363_/Y vssd1 vssd1 vccd1 vccd1 _2695_/Q sky130_fd_sc_hd__dfrtp_1
X_1577_ _1581_/B _1581_/C _1577_/C vssd1 vssd1 vccd1 vccd1 _1577_/X sky130_fd_sc_hd__and3_1
XFILLER_58_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2129_ _2130_/A _2130_/B vssd1 vssd1 vccd1 vccd1 _2129_/Y sky130_fd_sc_hd__nand2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2812__15 vssd1 vssd1 vccd1 vccd1 _2812__15/HI o_io_oeb[1] sky130_fd_sc_hd__conb_1
XFILLER_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1500_ _1504_/A _1519_/A _1499_/Y vssd1 vssd1 vccd1 vccd1 _1545_/A sky130_fd_sc_hd__a21o_1
X_2480_ _2481_/A vssd1 vssd1 vccd1 vccd1 _2480_/Y sky130_fd_sc_hd__inv_2
X_1431_ _1440_/A _1435_/A _1431_/C vssd1 vssd1 vccd1 vccd1 _1446_/B sky130_fd_sc_hd__and3_1
X_1362_ _2753_/Q _1362_/B vssd1 vssd1 vccd1 vccd1 _1406_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1629_ _1637_/A _1644_/A _1644_/B vssd1 vssd1 vccd1 vccd1 _1629_/X sky130_fd_sc_hd__or3_1
X_2678_ _2727_/CLK _2678_/D vssd1 vssd1 vccd1 vccd1 _2678_/Q sky130_fd_sc_hd__dfxtp_1
X_2747_ _2758_/CLK _2747_/D _2467_/Y vssd1 vssd1 vccd1 vccd1 _2747_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1980_ _1975_/Y _1977_/Y _1978_/Y _1979_/X vssd1 vssd1 vccd1 vccd1 _1992_/B sky130_fd_sc_hd__o211a_1
XFILLER_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2463_ _2463_/A vssd1 vssd1 vccd1 vccd1 _2463_/Y sky130_fd_sc_hd__inv_2
X_2601_ _2601_/A vssd1 vssd1 vccd1 vccd1 _2655_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2532_ _2527_/A _2525_/A _2521_/X _2577_/A vssd1 vssd1 vccd1 vccd1 _2533_/B sky130_fd_sc_hd__a31o_1
X_1414_ _1409_/Y _1411_/X _1420_/A vssd1 vssd1 vccd1 vccd1 _1414_/X sky130_fd_sc_hd__a21o_1
X_1345_ _2059_/A _1345_/B vssd1 vssd1 vccd1 vccd1 _1488_/B sky130_fd_sc_hd__xnor2_1
X_2394_ _2706_/Q _2393_/C _2707_/Q vssd1 vssd1 vccd1 vccd1 _2395_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1894_ _1894_/A _2728_/Q vssd1 vssd1 vccd1 vccd1 _2165_/A sky130_fd_sc_hd__and2_1
X_1963_ _1963_/A _1960_/C vssd1 vssd1 vccd1 vccd1 _1964_/B sky130_fd_sc_hd__or2b_1
X_2515_ _2784_/Q _2514_/A _2503_/A vssd1 vssd1 vccd1 vccd1 _2515_/Y sky130_fd_sc_hd__a21oi_1
X_2446_ _2470_/A vssd1 vssd1 vccd1 vccd1 _2451_/A sky130_fd_sc_hd__buf_2
X_2377_ _2701_/Q _2382_/C vssd1 vssd1 vccd1 vccd1 _2383_/B sky130_fd_sc_hd__and2_1
X_1328_ _2760_/Q _2692_/Q vssd1 vssd1 vccd1 vccd1 _1329_/A sky130_fd_sc_hd__and2_1
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2300_ _2300_/A _2307_/D vssd1 vssd1 vccd1 vccd1 _2672_/D sky130_fd_sc_hd__nor2_1
X_2231_ _2225_/B _2219_/A _2230_/X vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2093_ _2093_/A _2093_/B vssd1 vssd1 vccd1 vccd1 _2093_/X sky130_fd_sc_hd__or2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2162_ _2163_/A _2165_/A vssd1 vssd1 vccd1 vccd1 _2162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1946_ _1948_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1964_/A sky130_fd_sc_hd__xnor2_1
X_1877_ _1877_/A _1976_/A vssd1 vssd1 vccd1 vccd1 _1878_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2429_ _2721_/Q _2428_/C _2722_/Q vssd1 vssd1 vccd1 vccd1 _2430_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1800_ _1807_/B vssd1 vssd1 vccd1 vccd1 _1904_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1662_ _1901_/A _1661_/C _1661_/B vssd1 vssd1 vccd1 vccd1 _1662_/Y sky130_fd_sc_hd__a21oi_1
X_1731_ _1731_/A _1731_/B vssd1 vssd1 vccd1 vccd1 _1745_/A sky130_fd_sc_hd__xnor2_2
X_2780_ _2783_/CLK _2780_/D vssd1 vssd1 vccd1 vccd1 _2780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _1898_/B _1619_/C _1592_/B vssd1 vssd1 vccd1 vccd1 _1614_/B sky130_fd_sc_hd__a21o_1
X_2214_ _2221_/A _2216_/A vssd1 vssd1 vccd1 vccd1 _2215_/B sky130_fd_sc_hd__and2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2076_ _2146_/A vssd1 vssd1 vccd1 vccd1 _2099_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2818__21 vssd1 vssd1 vccd1 vccd1 _2818__21/HI o_io_oeb[7] sky130_fd_sc_hd__conb_1
X_2145_ _2149_/A _2053_/A _2154_/A _2054_/A vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__a31o_1
X_1929_ _1929_/A _1929_/B vssd1 vssd1 vccd1 vccd1 _1951_/A sky130_fd_sc_hd__xnor2_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2763_ _2793_/CLK _2763_/D _2486_/Y vssd1 vssd1 vccd1 vccd1 _2763_/Q sky130_fd_sc_hd__dfrtp_1
X_1576_ _1576_/A _1595_/A vssd1 vssd1 vccd1 vccd1 _1581_/C sky130_fd_sc_hd__and2_1
X_1645_ _1638_/B _1632_/X _1638_/A vssd1 vssd1 vccd1 vccd1 _1645_/Y sky130_fd_sc_hd__o21ai_1
X_1714_ _1714_/A _1739_/A vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__or2_1
X_2694_ _2802_/CLK _2694_/D _2362_/Y vssd1 vssd1 vccd1 vccd1 _2694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ _2059_/A _2121_/A _2121_/B vssd1 vssd1 vccd1 vccd1 _2117_/A sky130_fd_sc_hd__and3_1
X_2128_ _2113_/X _2126_/Y _2127_/X _2122_/X _2057_/A vssd1 vssd1 vccd1 vccd1 _2742_/D
+ sky130_fd_sc_hd__a32o_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1430_ _1430_/A _1430_/B vssd1 vssd1 vccd1 vccd1 _1431_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1361_ _2752_/Q _1410_/B _1410_/A vssd1 vssd1 vccd1 vccd1 _1362_/B sky130_fd_sc_hd__o21a_1
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2746_ _2758_/CLK _2746_/D _2466_/Y vssd1 vssd1 vccd1 vccd1 _2746_/Q sky130_fd_sc_hd__dfrtp_2
X_1559_ _1579_/B _1559_/B vssd1 vssd1 vccd1 vccd1 _1595_/A sky130_fd_sc_hd__xnor2_2
X_1628_ _1626_/Y _1624_/C _1630_/A vssd1 vssd1 vccd1 vccd1 _1644_/B sky130_fd_sc_hd__o21a_1
X_2677_ _2727_/CLK _2677_/D vssd1 vssd1 vccd1 vccd1 _2677_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2600_ _2600_/A _2600_/B vssd1 vssd1 vccd1 vccd1 _2601_/A sky130_fd_sc_hd__and2_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1413_ _1412_/Y _1412_/B _1413_/S vssd1 vssd1 vccd1 vccd1 _1420_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2462_ _2463_/A vssd1 vssd1 vccd1 vccd1 _2462_/Y sky130_fd_sc_hd__inv_2
X_2393_ _2707_/Q _2706_/Q _2393_/C vssd1 vssd1 vccd1 vccd1 _2397_/B sky130_fd_sc_hd__and3_1
X_2531_ _2577_/A _2773_/Q _2525_/A _2521_/X _2445_/A vssd1 vssd1 vccd1 vccd1 _2531_/X
+ sky130_fd_sc_hd__a41o_1
X_1344_ _2744_/Q _1341_/B _1512_/A vssd1 vssd1 vccd1 vccd1 _1345_/B sky130_fd_sc_hd__o21a_1
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_7_0_i_clk clkbuf_3_7_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_i_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_2729_ _2802_/CLK _2729_/D _2444_/Y vssd1 vssd1 vccd1 vccd1 _2729_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1962_ _1981_/A _1962_/B vssd1 vssd1 vccd1 vccd1 _1991_/A sky130_fd_sc_hd__and2_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1893_ _1894_/A vssd1 vssd1 vccd1 vccd1 _1893_/Y sky130_fd_sc_hd__inv_2
X_2376_ _2376_/A vssd1 vssd1 vccd1 vccd1 _2700_/D sky130_fd_sc_hd__clkbuf_1
X_2514_ _2514_/A _2514_/B vssd1 vssd1 vccd1 vccd1 _2783_/D sky130_fd_sc_hd__nor2_1
X_2445_ _2445_/A vssd1 vssd1 vccd1 vccd1 _2470_/A sky130_fd_sc_hd__buf_2
XFILLER_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1327_ _2760_/Q _1327_/B vssd1 vssd1 vccd1 vccd1 _2692_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2230_ _2215_/B _2225_/C _2218_/C _2227_/A vssd1 vssd1 vccd1 vccd1 _2230_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2092_ _2093_/A _2093_/B vssd1 vssd1 vccd1 vccd1 _2092_/Y sky130_fd_sc_hd__nand2_1
X_2161_ _2043_/X _2159_/Y _2160_/X _2146_/X _2731_/Q vssd1 vssd1 vccd1 vccd1 _2731_/D
+ sky130_fd_sc_hd__a32o_1
X_1945_ _1945_/A _1945_/B vssd1 vssd1 vccd1 vccd1 _1983_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1876_ _1876_/A vssd1 vssd1 vccd1 vccd1 _1976_/A sky130_fd_sc_hd__clkbuf_2
X_2428_ _2721_/Q _2722_/Q _2428_/C vssd1 vssd1 vccd1 vccd1 _2432_/B sky130_fd_sc_hd__and3_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2359_ _2445_/A vssd1 vssd1 vccd1 vccd1 _2503_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1592_ _1898_/B _1592_/B _1619_/C vssd1 vssd1 vccd1 vccd1 _1614_/A sky130_fd_sc_hd__nand3_1
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1661_ _1901_/A _1661_/B _1661_/C vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__and3_1
X_1730_ _1743_/A _1758_/A vssd1 vssd1 vccd1 vccd1 _1903_/A sky130_fd_sc_hd__nand2_2
XFILLER_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2213_ _2798_/Q _2199_/Y _2212_/X vssd1 vssd1 vccd1 vccd1 _2216_/A sky130_fd_sc_hd__a21oi_1
X_2144_ _2144_/A vssd1 vssd1 vccd1 vccd1 _2144_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2075_ _2075_/A _2079_/A vssd1 vssd1 vccd1 vccd1 _2075_/X sky130_fd_sc_hd__or2_1
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_6_0_i_clk clkbuf_4_7_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2802_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1859_ _1927_/A vssd1 vssd1 vccd1 vccd1 _1948_/A sky130_fd_sc_hd__clkbuf_2
X_1928_ _1928_/A _1935_/C vssd1 vssd1 vccd1 vccd1 _1929_/B sky130_fd_sc_hd__or2_1
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1713_ _1713_/A _1739_/A _1713_/C vssd1 vssd1 vccd1 vccd1 _1713_/X sky130_fd_sc_hd__or3_1
X_2762_ _2769_/CLK _2762_/D _2485_/Y vssd1 vssd1 vccd1 vccd1 _2762_/Q sky130_fd_sc_hd__dfrtp_1
X_1575_ _1898_/B _1592_/B vssd1 vssd1 vccd1 vccd1 _1619_/B sky130_fd_sc_hd__nand2_1
X_1644_ _1644_/A _1644_/B vssd1 vssd1 vccd1 vccd1 _1658_/A sky130_fd_sc_hd__or2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2693_ _2802_/CLK _2693_/D _2361_/Y vssd1 vssd1 vccd1 vccd1 _2693_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _2130_/A _2130_/B _2057_/A vssd1 vssd1 vccd1 vccd1 _2127_/X sky130_fd_sc_hd__a21o_1
X_2058_ _2058_/A _2126_/A vssd1 vssd1 vccd1 vccd1 _2121_/B sky130_fd_sc_hd__and2_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1360_ _1360_/A _1360_/B vssd1 vssd1 vccd1 vccd1 _1410_/B sky130_fd_sc_hd__or2_1
Xoutput2 _2199_/Y vssd1 vssd1 vccd1 vccd1 o_display_anode[0] sky130_fd_sc_hd__buf_2
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_i_clk clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2676_ _2760_/CLK _2676_/D vssd1 vssd1 vccd1 vccd1 _2676_/Q sky130_fd_sc_hd__dfxtp_1
X_2745_ _2758_/CLK _2745_/D _2465_/Y vssd1 vssd1 vccd1 vccd1 _2745_/Q sky130_fd_sc_hd__dfrtp_1
X_1558_ _1578_/A _1578_/B _1897_/C vssd1 vssd1 vccd1 vccd1 _1559_/B sky130_fd_sc_hd__a21o_1
X_1627_ _1624_/B _1624_/C _1626_/Y _1630_/A vssd1 vssd1 vccd1 vccd1 _1644_/A sky130_fd_sc_hd__a211oi_2
X_1489_ _1489_/A _1489_/B vssd1 vssd1 vccd1 vccd1 _1490_/A sky130_fd_sc_hd__and2_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_i_clk clkbuf_3_3_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2530_ _2590_/A vssd1 vssd1 vccd1 vccd1 _2577_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1412_ _1412_/A _1412_/B vssd1 vssd1 vccd1 vccd1 _1412_/Y sky130_fd_sc_hd__nand2_1
X_1343_ _2745_/Q vssd1 vssd1 vccd1 vccd1 _2059_/A sky130_fd_sc_hd__clkbuf_2
X_2392_ _2706_/Q _2393_/C vssd1 vssd1 vccd1 vccd1 _2706_/D sky130_fd_sc_hd__xor2_1
X_2461_ _2463_/A vssd1 vssd1 vccd1 vccd1 _2461_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2659_ _2673_/CLK _2659_/D vssd1 vssd1 vccd1 vccd1 _2659_/Q sky130_fd_sc_hd__dfxtp_1
X_2728_ _2802_/CLK _2728_/D _2443_/Y vssd1 vssd1 vccd1 vccd1 _2728_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1961_ _1965_/B _1960_/C _1965_/C vssd1 vssd1 vccd1 vccd1 _1962_/B sky130_fd_sc_hd__a21o_1
X_1892_ _1889_/X _1890_/Y _1891_/X _1883_/A vssd1 vssd1 vccd1 vccd1 _1892_/X sky130_fd_sc_hd__o2bb2a_1
X_2513_ _2783_/Q _2512_/B _2546_/A vssd1 vssd1 vccd1 vccd1 _2514_/B sky130_fd_sc_hd__o21ai_1
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2375_ _2380_/A _2375_/B _2375_/C vssd1 vssd1 vccd1 vccd1 _2376_/A sky130_fd_sc_hd__and3_1
X_1326_ _2694_/Q vssd1 vssd1 vccd1 vccd1 _1326_/Y sky130_fd_sc_hd__inv_2
X_2444_ _2444_/A vssd1 vssd1 vccd1 vccd1 _2444_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_i_clk clkbuf_2_1_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2160_ _2163_/A _1894_/A _2728_/Q _2731_/Q vssd1 vssd1 vccd1 vccd1 _2160_/X sky130_fd_sc_hd__a31o_1
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2091_ _2088_/X _2089_/Y _2090_/X _2077_/X _2064_/A vssd1 vssd1 vccd1 vccd1 _2754_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1944_ _1941_/A _1937_/X _1951_/A vssd1 vssd1 vccd1 vccd1 _1945_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1875_ _1875_/A _1890_/A vssd1 vssd1 vccd1 vccd1 _1879_/A sky130_fd_sc_hd__and2_1
X_2427_ _2721_/Q _2428_/C vssd1 vssd1 vccd1 vccd1 _2721_/D sky130_fd_sc_hd__xor2_1
Xclkbuf_4_2_0_i_clk clkbuf_4_3_0_i_clk/A vssd1 vssd1 vccd1 vccd1 _2788_/CLK sky130_fd_sc_hd__clkbuf_2
X_2289_ _2293_/C vssd1 vssd1 vccd1 vccd1 _2289_/Y sky130_fd_sc_hd__inv_2
X_2358_ _2636_/A vssd1 vssd1 vccd1 vccd1 _2358_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ _1591_/A _1591_/B vssd1 vssd1 vccd1 vccd1 _1612_/B sky130_fd_sc_hd__xnor2_1
X_1660_ _1901_/A _1661_/C vssd1 vssd1 vccd1 vccd1 _1680_/A sky130_fd_sc_hd__xnor2_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2802_/Q _2235_/A _2235_/B _2806_/Q vssd1 vssd1 vccd1 vccd1 _2212_/X sky130_fd_sc_hd__a22o_1
X_2143_ _2137_/X _2141_/Y _2142_/X _2122_/X _2142_/A vssd1 vssd1 vccd1 vccd1 _2737_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2074_ _2075_/A _2079_/A vssd1 vssd1 vccd1 vccd1 _2074_/Y sky130_fd_sc_hd__nand2_1
X_1927_ _1927_/A _1948_/B vssd1 vssd1 vccd1 vccd1 _1941_/A sky130_fd_sc_hd__or2_1
X_1858_ _1870_/A _1870_/B vssd1 vssd1 vccd1 vccd1 _1858_/X sky130_fd_sc_hd__and2_1
XFILLER_39_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1789_ _1789_/A _1789_/B vssd1 vssd1 vccd1 vccd1 _1920_/A sky130_fd_sc_hd__nor2_2
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1643_ _1643_/A _1643_/B vssd1 vssd1 vccd1 vccd1 _1643_/Y sky130_fd_sc_hd__xnor2_1
X_1712_ _1714_/A _1712_/B vssd1 vssd1 vccd1 vccd1 _1712_/Y sky130_fd_sc_hd__xnor2_1
X_2692_ _2802_/CLK _2692_/D _2358_/X vssd1 vssd1 vccd1 vccd1 _2692_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2761_ _2793_/CLK _2761_/D _2484_/Y vssd1 vssd1 vccd1 vccd1 _2761_/Q sky130_fd_sc_hd__dfrtp_1
X_1574_ _1898_/A _1577_/C vssd1 vssd1 vccd1 vccd1 _1592_/B sky130_fd_sc_hd__xor2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _2126_/A vssd1 vssd1 vccd1 vccd1 _2126_/Y sky130_fd_sc_hd__inv_2
X_2057_ _2057_/A _2130_/A _2130_/B vssd1 vssd1 vccd1 vccd1 _2126_/A sky130_fd_sc_hd__and3_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput3 _2235_/A vssd1 vssd1 vccd1 vccd1 o_display_anode[1] sky130_fd_sc_hd__buf_2
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1626_ _1899_/B _1626_/B vssd1 vssd1 vccd1 vccd1 _1626_/Y sky130_fd_sc_hd__nor2_1
X_2675_ _2760_/CLK _2675_/D vssd1 vssd1 vccd1 vccd1 _2675_/Q sky130_fd_sc_hd__dfxtp_1
X_2744_ _2758_/CLK _2744_/D _2463_/Y vssd1 vssd1 vccd1 vccd1 _2744_/Q sky130_fd_sc_hd__dfrtp_2
X_1557_ _1561_/A _1557_/B _1557_/C vssd1 vssd1 vccd1 vccd1 _1897_/C sky130_fd_sc_hd__and3_1
X_1488_ _1496_/B _1488_/B _1490_/B vssd1 vssd1 vccd1 vccd1 _1488_/X sky130_fd_sc_hd__and3b_1
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2109_ _2104_/X _2108_/Y _2104_/A _2086_/X vssd1 vssd1 vccd1 vccd1 _2748_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2460_ _2463_/A vssd1 vssd1 vccd1 vccd1 _2460_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1411_ _2752_/Q _1422_/B vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__xor2_1
X_1342_ _2744_/Q _1342_/B vssd1 vssd1 vccd1 vccd1 _1504_/A sky130_fd_sc_hd__xor2_1
X_2391_ _2393_/C _2391_/B vssd1 vssd1 vccd1 vccd1 _2705_/D sky130_fd_sc_hd__nor2_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1609_ _1619_/C _1586_/X _1587_/Y vssd1 vssd1 vccd1 vccd1 _1618_/A sky130_fd_sc_hd__a21o_1
X_2727_ _2727_/CLK _2727_/D vssd1 vssd1 vccd1 vccd1 _2727_/Q sky130_fd_sc_hd__dfxtp_1
X_2658_ _2691_/Q _2658_/D vssd1 vssd1 vccd1 vccd1 _2658_/Q sky130_fd_sc_hd__dfxtp_2
X_2589_ _2802_/Q _2632_/B _2588_/X _2183_/A vssd1 vssd1 vccd1 vccd1 _2590_/B sky130_fd_sc_hd__a22oi_2
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1960_ _1965_/B _1965_/C _1960_/C vssd1 vssd1 vccd1 vccd1 _1981_/A sky130_fd_sc_hd__nand3_1
X_1891_ _1879_/A _1985_/A _1879_/B vssd1 vssd1 vccd1 vccd1 _1891_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2512_ _2783_/Q _2512_/B vssd1 vssd1 vccd1 vccd1 _2514_/A sky130_fd_sc_hd__and2_1
X_2443_ _2444_/A vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2374_ _2382_/C vssd1 vssd1 vccd1 vccd1 _2375_/C sky130_fd_sc_hd__clkinv_2
X_1325_ _2771_/Q _1327_/B _2170_/A vssd1 vssd1 vccd1 vccd1 _2771_/D sky130_fd_sc_hd__a21o_1
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2090_ _2093_/A _2063_/A _2097_/A _2064_/A vssd1 vssd1 vccd1 vccd1 _2090_/X sky130_fd_sc_hd__a31o_1
XFILLER_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1943_ _1951_/B _1945_/A vssd1 vssd1 vccd1 vccd1 _1943_/X sky130_fd_sc_hd__xor2_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1874_ _1877_/A _1876_/A vssd1 vssd1 vccd1 vccd1 _1890_/A sky130_fd_sc_hd__xor2_2
X_2426_ _2428_/C _2426_/B vssd1 vssd1 vccd1 vccd1 _2720_/D sky130_fd_sc_hd__nor2_1
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2288_ _2668_/Q _2288_/B vssd1 vssd1 vccd1 vccd1 _2293_/C sky130_fd_sc_hd__and2_1
XFILLER_44_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2357_ _2691_/Q _2380_/A vssd1 vssd1 vccd1 vccd1 _2691_/D sky130_fd_sc_hd__xnor2_1
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _1590_/A _1590_/B vssd1 vssd1 vccd1 vccd1 _1612_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2073_ _2113_/A vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__clkbuf_2
X_2211_ _2799_/Q _2199_/Y _2210_/X vssd1 vssd1 vccd1 vccd1 _2221_/A sky130_fd_sc_hd__a21oi_2
X_2142_ _2142_/A _2144_/A vssd1 vssd1 vccd1 vccd1 _2142_/X sky130_fd_sc_hd__or2_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1926_ _1928_/A _1935_/C vssd1 vssd1 vccd1 vccd1 _1948_/B sky130_fd_sc_hd__xnor2_1
X_1857_ _1857_/A _1927_/A vssd1 vssd1 vccd1 vccd1 _1870_/A sky130_fd_sc_hd__xor2_2
X_1788_ _1793_/C _2001_/A _1793_/A vssd1 vssd1 vccd1 vccd1 _1789_/B sky130_fd_sc_hd__a21oi_1
X_2409_ _2411_/B _2409_/B vssd1 vssd1 vccd1 vccd1 _2713_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1642_ _1642_/A _1642_/B vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__nand2_1
X_2760_ _2760_/CLK _2760_/D vssd1 vssd1 vccd1 vccd1 _2760_/Q sky130_fd_sc_hd__dfxtp_1
X_1711_ _1711_/A _1711_/B vssd1 vssd1 vccd1 vccd1 _1712_/B sky130_fd_sc_hd__nand2_1
X_2691_ _2807_/CLK _2691_/D vssd1 vssd1 vccd1 vccd1 _2691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1573_ _1573_/A _1573_/B vssd1 vssd1 vccd1 vccd1 _1585_/A sky130_fd_sc_hd__xor2_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _2121_/B _2124_/Y _2058_/A _2086_/X vssd1 vssd1 vccd1 vccd1 _2743_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2056_ _2056_/A _2132_/A _2138_/A vssd1 vssd1 vccd1 vccd1 _2130_/B sky130_fd_sc_hd__and3_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1909_ _2006_/A _2005_/B _2030_/A vssd1 vssd1 vccd1 vccd1 _1909_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput4 _2235_/B vssd1 vssd1 vccd1 vccd1 o_display_anode[2] sky130_fd_sc_hd__buf_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2743_ _2758_/CLK _2743_/D _2462_/Y vssd1 vssd1 vccd1 vccd1 _2743_/Q sky130_fd_sc_hd__dfrtp_1
X_1556_ _1561_/A _1557_/B _1557_/C _1565_/C _1555_/Y vssd1 vssd1 vccd1 vccd1 _1578_/B
+ sky130_fd_sc_hd__a311o_2
X_1625_ _1899_/C _1641_/A _1641_/B vssd1 vssd1 vccd1 vccd1 _1638_/B sky130_fd_sc_hd__nor3_2
X_2674_ _2760_/CLK _2674_/D vssd1 vssd1 vccd1 vccd1 _2674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1487_ _1546_/A _1546_/B _1483_/A vssd1 vssd1 vccd1 vccd1 _1490_/B sky130_fd_sc_hd__a21o_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2108_ _2104_/A _2110_/A _2105_/X vssd1 vssd1 vccd1 vccd1 _2108_/Y sky130_fd_sc_hd__o21ai_1
X_2039_ _2054_/A _1510_/A _2055_/A _2142_/A vssd1 vssd1 vccd1 vccd1 _2039_/X sky130_fd_sc_hd__a211o_1
XFILLER_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1410_ _1410_/A _1410_/B vssd1 vssd1 vccd1 vccd1 _1422_/B sky130_fd_sc_hd__nand2_1
X_1341_ _1512_/A _1341_/B vssd1 vssd1 vccd1 vccd1 _1342_/B sky130_fd_sc_hd__nand2_1
X_2390_ _2705_/Q _2390_/B vssd1 vssd1 vccd1 vccd1 _2391_/B sky130_fd_sc_hd__nor2_1
X_2726_ _2726_/CLK _2726_/D vssd1 vssd1 vccd1 vccd1 _2726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1608_ _1608_/A _1608_/B vssd1 vssd1 vccd1 vccd1 _1630_/A sky130_fd_sc_hd__nand2_1
X_1539_ _1539_/A _1539_/B vssd1 vssd1 vccd1 vccd1 _1539_/X sky130_fd_sc_hd__and2_1
X_2657_ _2691_/Q _2657_/D vssd1 vssd1 vccd1 vccd1 _2657_/Q sky130_fd_sc_hd__dfxtp_2
X_2588_ _2798_/Q _2806_/Q _2787_/Q vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1890_ _1890_/A _1890_/B vssd1 vssd1 vccd1 vccd1 _1890_/Y sky130_fd_sc_hd__xnor2_1
X_2442_ _2727_/Q _2442_/B vssd1 vssd1 vccd1 vccd1 _2727_/D sky130_fd_sc_hd__xnor2_1
X_2373_ _2699_/Q _2700_/Q _2373_/C vssd1 vssd1 vccd1 vccd1 _2382_/C sky130_fd_sc_hd__and3_1
X_2511_ _2511_/A _2511_/B _2512_/B vssd1 vssd1 vccd1 vccd1 _2782_/D sky130_fd_sc_hd__nor3_1
XFILLER_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1324_ _2695_/Q vssd1 vssd1 vccd1 vccd1 _2170_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2709_ _2757_/CLK _2709_/D vssd1 vssd1 vccd1 vccd1 _2709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1942_ _1942_/A _2018_/A vssd1 vssd1 vccd1 vccd1 _1945_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1873_ _1866_/X _1869_/Y _1872_/X vssd1 vssd1 vccd1 vccd1 _1876_/A sky130_fd_sc_hd__o21ai_2
X_2425_ _2720_/Q _2425_/B vssd1 vssd1 vccd1 vccd1 _2426_/B sky130_fd_sc_hd__nor2_1
X_2356_ _2356_/A _2356_/B _2356_/C vssd1 vssd1 vccd1 vccd1 _2380_/A sky130_fd_sc_hd__or3_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2287_ _2288_/B _2287_/B vssd1 vssd1 vccd1 vccd1 _2667_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2803_/Q _2235_/A _2235_/B _2807_/Q vssd1 vssd1 vccd1 vccd1 _2210_/X sky130_fd_sc_hd__a22o_1
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2072_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2113_/A sky130_fd_sc_hd__clkbuf_2
X_2141_ _2142_/A _2144_/A vssd1 vssd1 vccd1 vccd1 _2141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1925_ _1936_/B vssd1 vssd1 vccd1 vccd1 _1925_/Y sky130_fd_sc_hd__inv_2
X_1856_ _1856_/A _1856_/B vssd1 vssd1 vccd1 vccd1 _1927_/A sky130_fd_sc_hd__or2_1
X_1787_ _1807_/B _1802_/A vssd1 vssd1 vccd1 vccd1 _1817_/B sky130_fd_sc_hd__or2_1
X_2339_ _2339_/A _2343_/B vssd1 vssd1 vccd1 vccd1 _2340_/A sky130_fd_sc_hd__and2_1
X_2408_ _2712_/Q _2407_/C _2713_/Q vssd1 vssd1 vccd1 vccd1 _2409_/B sky130_fd_sc_hd__a21oi_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2690_ _2727_/CLK _2690_/D vssd1 vssd1 vccd1 vccd1 _2690_/Q sky130_fd_sc_hd__dfxtp_1
X_1572_ _1898_/A _1577_/C vssd1 vssd1 vccd1 vccd1 _1573_/B sky130_fd_sc_hd__nand2_1
X_1641_ _1641_/A _1641_/B vssd1 vssd1 vccd1 vccd1 _1643_/A sky130_fd_sc_hd__or2_1
X_1710_ _1710_/A _1710_/B vssd1 vssd1 vccd1 vccd1 _1734_/B sky130_fd_sc_hd__xor2_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _2058_/A _2126_/A _2105_/X vssd1 vssd1 vccd1 vccd1 _2124_/Y sky130_fd_sc_hd__o21ai_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2055_ _2055_/A _2055_/B _2144_/A vssd1 vssd1 vccd1 vccd1 _2138_/A sky130_fd_sc_hd__and3_1
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1908_ _1995_/A vssd1 vssd1 vccd1 vccd1 _2030_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1839_ _2735_/Q _1839_/B vssd1 vssd1 vccd1 vccd1 _1851_/A sky130_fd_sc_hd__xnor2_2
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput5 _2234_/Y vssd1 vssd1 vccd1 vccd1 o_display_anode[3] sky130_fd_sc_hd__buf_2
XFILLER_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2742_ _2759_/CLK _2742_/D _2461_/Y vssd1 vssd1 vccd1 vccd1 _2742_/Q sky130_fd_sc_hd__dfrtp_1
X_1555_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1555_/Y sky130_fd_sc_hd__inv_2
X_1624_ _1899_/B _1624_/B _1624_/C vssd1 vssd1 vccd1 vccd1 _1641_/B sky130_fd_sc_hd__and3_1
X_2673_ _2673_/CLK _2673_/D vssd1 vssd1 vccd1 vccd1 _2673_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _1489_/A _1489_/B _1349_/A _1479_/A _1479_/B vssd1 vssd1 vccd1 vccd1 _1546_/A
+ sky130_fd_sc_hd__a311o_1
X_2107_ _2102_/B _2106_/Y _2749_/Q _2086_/X vssd1 vssd1 vccd1 vccd1 _2749_/D sky130_fd_sc_hd__a2bb2o_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _2055_/B vssd1 vssd1 vccd1 vccd1 _2142_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ _1360_/A vssd1 vssd1 vccd1 vccd1 _1341_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2725_ _2727_/CLK _2725_/D vssd1 vssd1 vccd1 vccd1 _2725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2656_ _2625_/X _2654_/X _2655_/X _2636_/X vssd1 vssd1 vccd1 vccd1 _2809_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1607_ _1606_/X _1599_/X _1899_/A _1612_/B vssd1 vssd1 vccd1 vccd1 _1608_/B sky130_fd_sc_hd__a211o_1
X_1469_ _1590_/A _1590_/B _1470_/A vssd1 vssd1 vccd1 vccd1 _1471_/A sky130_fd_sc_hd__o21ai_1
X_1538_ _1539_/B _1538_/B vssd1 vssd1 vccd1 vccd1 _1538_/Y sky130_fd_sc_hd__xnor2_1
X_2587_ _2587_/A vssd1 vssd1 vccd1 vccd1 _2587_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2510_ _2782_/Q _2781_/Q _2510_/C vssd1 vssd1 vccd1 vccd1 _2512_/B sky130_fd_sc_hd__and3_1
X_2441_ _2441_/A vssd1 vssd1 vccd1 vccd1 _2726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2372_ _2699_/Q _2373_/C _2700_/Q vssd1 vssd1 vccd1 vccd1 _2375_/B sky130_fd_sc_hd__a21o_1
X_1323_ _2692_/Q vssd1 vssd1 vccd1 vccd1 _1327_/B sky130_fd_sc_hd__inv_2
XFILLER_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2708_ _2807_/CLK _2708_/D vssd1 vssd1 vccd1 vccd1 _2708_/Q sky130_fd_sc_hd__dfxtp_1
X_2639_ _2805_/Q _2632_/Y _2638_/Y _2622_/C vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1941_ _1941_/A _1951_/A vssd1 vssd1 vccd1 vccd1 _1942_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1872_ _1871_/A _1871_/Y _1872_/S vssd1 vssd1 vccd1 vccd1 _1872_/X sky130_fd_sc_hd__mux2_1
X_2286_ _2667_/Q _2283_/A _2482_/B vssd1 vssd1 vccd1 vccd1 _2287_/B sky130_fd_sc_hd__o21ai_1
X_2424_ _2720_/Q _2425_/B vssd1 vssd1 vccd1 vccd1 _2428_/C sky130_fd_sc_hd__and2_1
X_2355_ _2355_/A _2355_/B _2355_/C _2355_/D vssd1 vssd1 vccd1 vccd1 _2356_/C sky130_fd_sc_hd__or4_1
XFILLER_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _2137_/X _2138_/Y _2139_/X _2122_/X _2055_/A vssd1 vssd1 vccd1 vccd1 _2738_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2071_ _2075_/A _2043_/X _2079_/A _2070_/X _2041_/A vssd1 vssd1 vccd1 vccd1 _2759_/D
+ sky130_fd_sc_hd__a32o_1
X_1924_ _1924_/A vssd1 vssd1 vccd1 vccd1 _1936_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1855_ _1854_/A _1847_/B _1854_/Y vssd1 vssd1 vccd1 vccd1 _1856_/B sky130_fd_sc_hd__a21o_1
X_1786_ _1786_/A _1793_/D vssd1 vssd1 vccd1 vccd1 _1802_/A sky130_fd_sc_hd__xnor2_2
X_2338_ _2688_/Q _2342_/C vssd1 vssd1 vccd1 vccd1 _2343_/B sky130_fd_sc_hd__nand2_1
X_2269_ _2666_/Q _2665_/Q _2668_/Q _2667_/Q vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__and4b_1
XFILLER_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2407_ _2713_/Q _2712_/Q _2407_/C vssd1 vssd1 vccd1 vccd1 _2411_/B sky130_fd_sc_hd__and3_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2815__18 vssd1 vssd1 vccd1 vccd1 _2815__18/HI o_io_oeb[4] sky130_fd_sc_hd__conb_1
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1640_ _1638_/A _1638_/B _1629_/X _1637_/Y _1639_/X vssd1 vssd1 vccd1 vccd1 _1640_/X
+ sky130_fd_sc_hd__o32a_2
X_1571_ _1571_/A _1571_/B vssd1 vssd1 vccd1 vccd1 _1898_/A sky130_fd_sc_hd__and2_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _2113_/X _2120_/Y _2121_/X _2122_/X _2121_/A vssd1 vssd1 vccd1 vccd1 _2744_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2054_ _2054_/A _2149_/A _2149_/B vssd1 vssd1 vccd1 vccd1 _2144_/A sky130_fd_sc_hd__and3_1
X_1907_ _1892_/X _1906_/X _2041_/A vssd1 vssd1 vccd1 vccd1 _1995_/A sky130_fd_sc_hd__a21bo_1
X_1838_ _2734_/Q _2733_/Q _2052_/B _1829_/B _1823_/A vssd1 vssd1 vccd1 vccd1 _1839_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1769_ _1792_/A _1793_/A _1793_/B _1793_/C _1768_/Y vssd1 vssd1 vccd1 vccd1 _1793_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput6 _2228_/A vssd1 vssd1 vccd1 vccd1 o_display_cathode[0] sky130_fd_sc_hd__buf_2
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2672_ _2673_/CLK _2672_/D vssd1 vssd1 vccd1 vccd1 _2672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2741_ _2759_/CLK _2741_/D _2460_/Y vssd1 vssd1 vccd1 vccd1 _2741_/Q sky130_fd_sc_hd__dfrtp_1
X_1554_ _1581_/A _1579_/B vssd1 vssd1 vccd1 vccd1 _1565_/C sky130_fd_sc_hd__nand2_1
X_1623_ _1626_/B _1641_/A vssd1 vssd1 vccd1 vccd1 _1638_/A sky130_fd_sc_hd__xnor2_2
X_1485_ _1485_/A _1485_/B _1485_/C vssd1 vssd1 vccd1 vccd1 _1489_/B sky130_fd_sc_hd__nand3_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

